XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���]2��J�����^�C�b���vw�˝nE�F�g4�C5ʀ�� 1�Lg�zuP�5T��8��s=�"c'I�a�[Hd?G�u��ě�T61�FɎ,�ќ5����_3A
u�j���߲V��x_R|��K�H�C��b.���Q�²dj29w�9q-�RX�y�r'sj��VK����^h Bh���a�U����������I�2�gƿ`�@��fQ}Ws�Ǒ;�U%)J$ǹ�����+Y8e�b�lH�/�;���=�vġ6\�G7@�vy��r�o�O1!K^���e����k����y��,��,Ԧs��Ѿc���pY���t>^TSj|[��7���vI�?��m��S�Sf\=0.����0�	�����]�K9+�9������5姗���j���L��>  4�;h�4%�-J%4��}X�8�`p���қb���l�et��#�<�K��z�����L�E9)y�ۓۜj����AZGO?	�#\��f���ʗ��_�x�/D��kPc�,��J���in
kmg������z���U��
�H�j��2<�~n�7*f[뵄���󺜍n~B��#G��C{��p��C+{e:�Y�-f,��-�_����'SP�\~���{'X�J�U���h@u�(�g5��c�O���`^�민Ӛ�D5e��k�88��et��=��Ǡ���s�n�4�F(T������^�z�5����&����,~9�B�֦XlxVHYEB    136d     800̝�G/.�x�&���jmh�a��:W����h�3���gc�󾥼��ْ	��M�������uZ����#M�é]��f�oA�C�+U�J_��?I�]#-3�f!R�����QA��5���J�ȁ<�{i�s��ip�|/�v�s>m�O2X>�F��R���:�S%Ն��l�q2�z�.e��~�ݚ�R4�Q���J��>����2���)8��- &Tփ�uԁhQ`l����� ʬF'u8,�(��z1\x�p��T:�hџ~�@��E�`x� �R�D���I�tO�х����k}0���G��r>�����>b>�ܛt=z.m�P�ofr4���U�w�i���s4X[���Y��m	o�j�ڲ`oӑ)BiƩ>!��̸�]X�б�AW�@o:	�Ź�8lp�c8^)������_��h�Q�/��RG��9*�(�����Mvs�v���4�zB9y�W��taz�qcSk�5���>z,�f��i�G�$.I���R%({�#H���>NC�O��%LS�>��O���_E@����V
ȗ�r|��Aȃ���Ŗ)�Y%�ܘ�m�q̠�K���S<��HG�;0k����A@n�O���A��`\�g���'����n{;u����(j �yt�P��(?$�
�d�B{[�w�ު�u�<	\%#_������������&D�u�7��2F���ec�DC�W&Ϙσ��}���2�OLNmQ[�x�%_�
4yO�D���2
���B�7h Ϣ�i�uh�v,f0sJ�RӨzNw�.��7��xyJR�%�^3������"�\������/&4'_���u��"��Z��"Gws���5p�RnNnD\��~j�� {��Rڤ<j;��X�nRV���\�-ˠ�o"O�|"�M�.�m
��5P��E7����g�ȡ��1��tz��K�4��/m����&E��Ղh~3�
���ň�=u�AF�D�dxT!J!��%���ZuB:7S �@�#�g.�t@����PGp��Ru�
o�X}������Aƺ�$4�x���0�ʐ]_l=��1�$�b���0u�<�369A��Tx�\2��b�9�2.�'K_,�n�`�o��q�#���I��PM4����O	
�J��Ӎ��B�W1p���� dd*�A m�_�qt[��=S���xbPX_	��9��K�w/B�[�	ւiƲBfR]���e����@N�;�2!7���Rvb�C�5Mϲ��o-�q��<��;��!���8W�}��4ik�)~R�����@�'L�׉��=�X�v���7wahT�64-a�%涽�2_��VA8b�Ϭ��Вt�kt��?`>����'0�C�E��x���/f~�� P}˳Y�YGc�t<�s� c�pH��3Z4ӗ��	G?�E%�ڻ���'���;07W�%�wj�d����Q�)o�>���W_מ4��	��TK�غQ G�FxF��y��t���S��3�GQ�A�p�K���2#"�rH�L.):�[p^�M�	*U$6&wNd �+�6��K�T�<����{��& �Ny�)St>�]����(O���ᷨ�P�io���F������='�݆��8"l�h=+��\(E5f#���ET����[��@U	H	�%p�R
��n0��R��!Fr��̹�#y^�$�j�,��٬=��v�[���0����V�p�E��H�:�K��� r&& �;9�x�e��Q��゛��@��x���Ҡ_��`���5>��j����+.�Eq�fn�8.2Z�d�۽wr���bgJ��l�(��]��Mr
@�㈺��!�4µ3f��r�-��U}����6ښ��o��	��=!es�י��+	�cU%X>ڦFnv�����;C�Lpŝ�\ºu��\I�i�����c�1v�=�up���=5#aj�z�Q
�_�T#�V�!�C�x�tԈ�rȫ�(Qw��ߣa�`�ڭgH���j2'U�`���a ɡ����4)��_��`B�;�0f��Ȇ