XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��������� �Λ�r�H�ϡ��v�v����K�QJ��q�dS��~Ӷ���u~	T���χ[����d
Y,_)��,_��0�<���j�)>w�?��`L .`�<�Df�Wi�~n@B�s���L�2�������>��f8&a~{&,:&��A��;1{��%����܁�__�-��_��.�M<[�l�� �io3&y�״`��U���HR��:i��9YL���j��岭6�mv���kw �z��gyJ�E;e�v�x�4���4��"��6�R�C�Av���8%�Dz<��I�[^���t�hGG�Ra�H�+8 yM�ó|r�t��+�K�)�\P��ۗ�gWZ�ROa'���ˡ ��:8F�p9Q67̒��r\��������0�]b�&�� m�u�]�*��\Z�amb&�08��&��_��K��l���~o@���E�SJ˱���@+#δ��8�P8�6� :�%�mW������l-uJ��������s0����jn�U��7#ϙ��[�Oy���r�XP|{�������yt4��yכ�� �W���+�hY���`Zv�&�{ơ��ϛ~\�b��"6hi�.��
r�Vt��F���ׁ��0�n�]n�#| ͬ�؆ϧ�M�
Qa>V��(��hA�L��Q@��8p�~��у��k��.��i��_
z�2L�2����	�N�4���T4��)��T���ޛ>�WW�l�i��F������CҐD��1d��� ��~��nRXlxVHYEB    eee5    2920q݄C���S�2�Gsqc!Ȉ�1&[���s�m����k��,A�/alB�YVy 6���1}[���x�d0��+���(����,���� ��1T�(:�{�!jP�+�:!��Ϩ�2��"���LO���v`Q�^8�0o�ګ�>�A�$dzOέ� +�|؉��}�dQ�0Qӄ�
��<G
���1�x\�l/�-؝����BIz6O��0P���<��C�#�׋WI�� ���z���K9G��z�=�j�qH[5�S��H�Ĳf�|<��{����V�>º�/v`���嗲|_ŏ�0�>z��A��#���N(@��赁T�sd��^y�($�� ������&�	D�Ս�a��U@V$��F���~�v���%�	X~�Œ�p��u ���lPj�]	~S,ɏ�ˈl�i�bdHM��LU���fEt�(�eۜ9Ogg5~sB9�X�K�G?�������Q'/����C�ʛ��~2H6�{�4�'�5?���h��w���u�s�}g���Te�_��l�-yd�`R��Q�b)o���U2=��B��	�d��YF_CfN�=���7�O��S3�g�'
�3�,:"�u_@dǲF�@��!-1WGg��@�r�ʀZ��=G�mW��K$�V 2�!Ԧ��8|�P$<���I���1�S�ڜ~���t{/z�y[��7]�e/��x⯷�ƚ��1qnR�U�X��Ąr����Y����ǚ�fҹ��rC���ԍ���H/%$[��3A<�j��B���4�`�k_>r�6}�1b��TW�4�v���gXl���T��]4J�~�3,I�B���B1�SWs��B`o��;2�ڀ4��oD�o&8�?39���	���9�Qy���W�����=����YPh���7&,
㸀�<�SU�E9��Uj��[��g���/����{������U`r�P�sZNr���<��J.5�y��EE���*�,���7ݡ$�>|��!����[u���5�g.J��a	�)�=�('�!oÄ�*]���{3.�Y�U�����*{a��\�76�-Nz�H?[�E�3b�&���o��"a"�"2���c�D��ez�*�|4햛�f���	'!�D������/��v�Ί��	�M3K!_�_�u�Z<��U��[e��fi�u��w	�ba�:��pg��Z_��g�EeE,�aD�r�2I��#�6�x7Kԏb��a|��u�'��T��LwhGP\���s̓����4��%8&#)V���ڝ�|��x� 4����7ػ�9�	8-x�HPD)���{�0[�qq~��'����i0o,��);!�צ�>�yO���R���g�z�P�q�oaKR;MK���*��#1���*F�NJ�\��}0���d�����4I3����3s>��*%�E։��y���χ*T`F��z�����͗'��8��v��9��F��7��L]�H�g��O��k�����p;��嫹Mx6F������^<�#m�\=,�%�������r���0�Iv��X�%�,&k���z�aw��ş�� UA��j6ck�Fg�1�+<֋R�t�hs:�l����C�������;�_����Z3��ɇBC��#����i�n��͹6���z>������\kk��uo��3O�����*��]��.�Z�4&"�ZXyt�0��A�Lm�݇�{1���'fU�X�e�m�i��Q5G�+B"$��=1�[�|C����M`��P�ޙe����2_B	}��hf�xz��zDS�O�7�hf��-xwf S�a�q��mvH#�"y9���E��P�F�I�O��ZĹ��>�T�\l<}\������K�DD�˾�:�YP���;�K-M������C��p"�ҥ`Ny��o'g����Ǒ�q̽\L%t,��h}5���jI�����Ħd���%�gSeY���΍�nU�ԤJq<3 �O�
��yk}����e�	,-��� 9����m>�� ϙt�ť��;QF�zD��Z�}{�+79�2�Aa4BSW�#$��%��=�/�׷����K��t`���1���Xm�R���}`&Ԥ��?� �đLF<EO������֛d�j�a�L���x�� Rm���sr8�������80����Ez�y���n��4�aj}��K��N8T'u0l>i	m�b�=v�@��W��AO��4#�Wp�*��l�S�|<�i�̌�;��c��Bl�Uu=�R�/s ?���)n=ƲM�W�27��w)M˚'�so���1������/�g%B@fgpW�~*�;�]~{��Ќ"z�z�T��U[g_c�,+��G���
v��%v1�[S��(;E/o\:e�'���λ��+a�����`߼
��)�2�?���JO��D!è���tB�l���pܫT �U'���Io��P��r��o\n ՄaL銻��%]����[�B��1AL"R�F5�'6�����9����CD������E�6,j)�`�O5Jj@k9�B�/8�haa�Y��{ɂ���v�( �٪H�� a��`H�O(�>O�� ��V2A�ٸ1	�
7�!�BQr�	-ʶ�.ͧF����Mѩ�����DᲃG[.t���P0D�6K�E}�(���)��s$Ly>��u���]��o}nlO�-X�w��Tп����ϤGJiS�BG�D=E���F�<�t��h �M=u�e;�M\2��O���d���Q|��x�5"���C:j�[���6j�X_� W-�����E���V���1+c�,R�߆kxbzPi�hC/��B�h�ud���k{�R�t�z����(P�V�jߞ5S��$b
�f P�R��	�a�(Q� j�3}?AY��+��,��H���a+�w��Ys�u(D��IZ4_5Sv��\����
����̿����	��#��:��K1B�0,��a�C;!�l���3^���>�(bY�/dG�Ⱦ��$ji��01��z�9�M���D~���o������Y@��L"���x�g�.j�Y��	���'��bR�$c�eb+M��Wag�[n��"}�2�/��nk�g|�\;c,gp&��Z������%�=�W��UbQ3Ïy��m��3v����^D#�ĴͶ�{R%J(|�J���C_害�V����]\"���S�r����O�D����h��f�+:�D�����L�O��������:H�%r�I���x4*f�%d��&�l32�F�1H�>n�d3�YI	�٩��k��k�emz��Ȍۄ܈R?�| ��`�>��72*�Q���ʜ����������r�1�G�����xc��w����g�ݺvzJw�n�&<��#(������_}JR]�0�^�k�_'�� F�y��8�B��q�2/��%x����x��t3|&Y �U���v����.j8���W����&X�0z/h�R��m-oUVg��qI��,5��K%��҂#ίbFzi�?�)%�Y%k�T!f HH^ոH7���q�_����t�HL�򻇄�P�ꋱ :p �a�OJ[���!����TreyN	�5Q-%���ΎJl#*Q���|VQ���Dvj��-gI5����Ơ~��(Ŭ�33�~�i�|&��d���v���/�Ջ]��C�9��۹�D-IB��/
��4��Nf�6,ɧ���Y����Э�fewٰ�쐞����sS�dꇉ��@����>G���|��Oh{��3`�;1꓃=iv��� ����xG�۪�ҋ�Ö�%�iy��[��w6\I��,M�l�׏hW��mκ�W\`�\�ڣ�jm��Gֳ4�ͼ#:7I3���h�CzV�k������5���z��gL1(��쏮��`vή���$�lH�\ѹE��2��p�$��/���D�3��v�����I뾺q���I��M<�ѷ�zpmv�)��4�x�sѭ%��-Ț�I�@�>7�[Y��������F(Nl��c>�H��Xp2T�b���U�&�M�L�����!YWK�<�܋Mv��׶ϗg�r�a�`6C����]�6}��6b������(u�qnAV;��T�Yi^�Q�d��:�x���%Ry�ᦐ�T4�W���`'ؙ�0�Z����ܵ|�U�3|�e��N�"��ɽ�c� ��"�B�������VrN���!̽O�>��fB��B'@��n4 �Zix�;Y��<?ւc�?[P�	���\��i����_����M�txC��y��ǭr�:]) ��g��$ԝ�Θ�`�Cο�St�dv2҅�Pa�Go����[ �n_b(�^k�N�W-�f��ٺ�;d�@��-����'9��R�V�J��en�������NFFJq�5r�b�t6a~�k��4ЃLgV�'�.��l�7�*��_gw�Njk-�-Sl��l].e���c7����Q�JD����|�ؿ��9	u柑�"$� g�j�B��MI��F�n� �"������Սr��<���
�
ٜž=���,��"����^���H��o�*Uc�.T�uX=�h�a�,��=�Fp�'�ّ�4FGǴ	a�9����4�2�.�  ��KG�1�i��S���?e�۾@2�0�"�z(M�$~Qj���kp5^�]�2juh�W���ć� ��m@e�@=���'��5����}v&��7d��X�������	���Q�t�ਓlaBGQ4��S��h��V�k?���P��c=���GJ+� 0�6���,��7'V���Td}���r�WA~-���*��5v��z���-|�ď?�bM���p�����LQ�訣T�:?}̛F�E�*b�CC��`B��$�
0�� �ոV�Q���l���{�ʏ?U�JS�����nܹ�(,1��Ǆ<+�d&�{���B���EBA��Q�@5h�E�)G�v9�7�aM��<�+�m�f� i/���H�"n(��}1T������{^4E����HR��f��:�J���F�Ȼ�r�#�6|NWa)!"�Ir�`,h�rx��J��7��L���pێ�;��*G����J�އs��}^���0x4�����G�ф��S��"p>o��!L��`�7Z���ʯ��}_q��,0e�@�?��l��9��kݍ;�[�`�z�����h��y&9�$�MB8*����l�C�'��x����~�ͱ1��:�3,�1��������=VEU@��n¬��EJ<k�P�G���h�Wi�G1ܨ#��;�i&@�߹����wmƗu���|P��\�Ķw��hbP"�X?�&��p@�c���?1���ǜʼ����+�7UC��xv��N/s�e���q0��sS�;�|`�`����g©�!<"g�W�n�6r���6Zn���(�J��w�(X��
��,�pAVd�g��Mv���z&���]��_�L*V��N���_��Z���k"6
<d�/�%#d�ҸHO�h���?J�,}�}t�������̍r������������ϒԊ�ÂVw΢��B���t��Í���&\�2�J�قcV�� ��{��.�i7GW���x���U��.Lt\���X6��]5��/v�<7)*l	d�5y�����r[�8F_�:z������_:<G����+.�Y��g���r1]��$s���P�-ME�jr��z���!|��G�{�S���ܑA����k���!:v|�zҞ;xD�#�����+pO��(�	-^�p�y����)g���̺n���&1�pckK���@��
��Ij��X�5�����Zj}� S"0Y�<oP��4�n�ټ"��!�90P E�Ϻ���I��"Wo��RN�k6�є�����-Zʗ�� ��[9����p�cZ�&$=��J�|!���lk��@�n�=_g,�Y�'����m{"ڏR8�"��0(�NXC ��!��ؑ(!r $w���m�����s�������鼈H+=#�J)څ|7�$�ڎ�S��C`�o��$d2���&~De��DKkm$��n���e�J��)e�ȍ�n�x��CM�`9��*O���㈖JV��g$k%y`)*�Q{��!���=g�zܺg ���E�S���s5(�
���u��6M{��l�7N������g<���H�_��g�>wP�!�.p�9K�u�n{̘����e1��I��m�ض�MCAE
�:�z�������\Ob����a�Xb-4@�(�O�>;�,�~�3�K{�$�\X w�n �� 3�[e(���6����W�0zJB=pj�P�jq����OԴ�2(�|��z�y�ȴ�Rӫ@p't=���ͶR"�0i �g0�3�]�hm�����l|Wn��j�O���*��[�s�ӷ��*��	Mz�(,���,�},���F`�gU�,2襜YN�3j�?�T�����.'
�1?R�PT�A�Q58V���P���&,Y�j��L��A�6�QW#�O�s�Һ	ݢ	�@�.�������ף�c�{�S*��W�W�.�����u���y����eq�U��:��U,�t����6�6�J�m�v,�n!�!T��'f �_!�#ܒS�X�ǝE�H�yJ�d�h�ӣ�m�6ȩ�h9J���~V��?�f�� {jH������4��3x�yE� _��b���4�]��^���2;XX.�ߚѯCO����Yo�4��ICir��Y_n�\�I*�]1ʬ��w2�)]�=�`:����6��aS���s�=���]l���+ed�Z�s�+/�)ڷ���BE�!P��sF.49�4��b�� [�i܅�]��^J���n�� ����!B��~y�ag��:h.B������)��Uդ�Z�ݝ,���K����$���:�X�>j u|�}&��-�W���I?~��s�K�+s�,�m����p��P��r��#'������u��.{�����%��`��)�b���:,�q�)L��y�"]��
�$J`�J��پ�(o���[�ZO�,l곛��?4'�6���IS�<������`������c�}� ��>�.{o����s��1߉�}�8�}��#�amY���Yd>��&�FKq�n���T���r�dz���S�ғq��]ݽtq[��N&Utz��٤0G�Vѩ�S=)�8�#E7q��ɋ�`���_*��Xp�S��f1Dp�l<�21��C�
4t-����E��F��\4YjpK�@r�����A�PJe+������C
I���F2��ڴ�H����a�(�1�[��6Ɓ�c
:���nj�(�2`�J�VMC�<J�I�56W�( �b�9���*ЋS���"��9-��o�sW�9�N�]OHP�]K���$�oжt@���AC��Em?@��w*P&�(�׮K�xs�/E>�r<m6�E�Z�h/2�"C��A
N�n>���]�"��}[`�A�l�r��V:��3�=Ø8`��0%��G=� ԓe; �X}|3*�2.��z�z�
��}gF1�fdD��#L���PE|�9�F�G��pw�"��3��w�m�32��5�$2�`~�����I��$Y˿�0Q��Ct'�Ά/�zN'͜�}`�J�m�rUkOQ��� �����CB�*��P���b�2�c�{pY�뤪��)�I��a���a�,6D�>{�n�IH��a���͇T?N?֒N1(ķt1 ��[��{؋-���oXwZ�������oT�i=iP�|�>��O��+�/B=`#�}�yz�o�V��?����n�3��B��z$���@$�$VȎo�n��z�=��!�ˤ�q�jB#r\,}e���9B��f��ΐ��$Rn��=7)r��Gu�^�M�O�b9q�٣����&�K]���I(�sJ�x:Z'� ��"�4�u�.�����\o�k`H^ @��"�n=��P�Uri�1�$u��_���� �d��F��e�rH9�"�zx?���A�6�8o*'d���Ƕ7�R���_�E�T�b�g�)v�A���dA��	2�8[X�"��f���P�G��ؙ��#����ȉ�s|�Ȕ\�H�g!F��<w���jZ�
;�F��E�%�O�0.����a>/-x�����ƃ1��7?��qX+:��v1K~o�mt۟�%��?�S�jE�v-��k.pFK����K�Jʅ��7j�r���o*���B�r�,#e��@�I�~p��$Iªͧ��3Q�C?�*�^>�����&hU_�p�&�[���Ï�ȕ<5��y $���>f;<6
`F�.A����ױ�UN�ϹQ�#�-���p�h�.\)� �E�FEDy���{Jᡅ�����^��A��v��(��i�\q�������N��7�-|K���[L�EM�9�yұ�?�>�����K�	�>ߚZ���(NV�엋}#�Kۏ�o)@3"�F�:>m6��i>^?f,��6����X��FѝmkR
Z����aVJ7�Nh��$1�.�HD'�n5t����1�R�[{*F|��]��eF�ݎ��K�<C�!o��+`��+�Bz�LH,{�6I��A����Gy��p�;6~~��jh�f��V�hl�FIm�~�=��Z ��@��\��>��Lm�HE/�?�{nQ̜�ť�C�O}�1�|����`d�M�i��\fa�!�X��b�ƊQ�#SK&�*QR�Gz �qNҲ���<r�>�[�aç&G�-ytM�h(�����3	�&��9@�]/d{�]~㢺b�u>%e���x����LIInI�4c������L"b1�O��p =zc�g*{� ���8"��1
sm6W�фέ�!�k^��B���DJ?M�Yl:�#�e��B�I�n|�_aoW|�Y��=o�����++���/���G1Tc�=���]��/�]ݏR��3���J��\<$�=d8<k�>�:	�^��M���P8������S�5����nV$j����?&�|�w�����Iz�_��z6F��C��]Fy1�+ؽs-��I\ܛ���y
���p�P���7�xJ�!L��M[\�$ݦh�����qR]�k�����$��#����,�I�$�'Nc�d���z�|�Y�C�ҌB"L�������r�ա��xn0<��Q~U�&����6�q�����R���g9��j��a��]��'�&ö�K���t���|��u� oXA?��)�lZ"�79�U��9�w�kYnOA��$�!�������M�И�F��"��s��oD"��7��R�}�|���� ���(R]$��u+�\�Qu:iIl������$����*.d����|�?�x�M7�
Rv������3��� ����Q���98'���u(,Pf!��9�i�p�7)5�d���.Q�q��\o����ft4e>�o�A�������	�zo����y����O,H����i���lǥ6$��d,�ΫUZR?���K��_�z�t�?��$)C����${�^��L�Z�4�����VK�&�r���]l�v�+ ���n A�v�K�8pYc���X?@�}�\�K�)����K��?�rG���2N�~�ۻ��]cF�>��w�]۶T�h�),����č_����㧔Y�!;���P)����r�b�h���'�h��8Z����������~�#����g?�#��Ohף��1���*�p�N�s�(�R�w��X%�>���c;�P��[=�� Pۅ�Ì�����ĩ���u:����B#����[I���(ώ|�l�{
� ��ǯ�:7�?�k;J4�~���+�㫞 tsT��Ȼ�د� N���"�����C�c�`fyìPZw5�P��f���H���M�3�W�q�by�\�$d�MO�.5�НL�Sk����/�\����?�Fj1Y�^�$�'k-�r?9�&,Pct���-AƷ��ԶE��Sz�.�i��G��~6d���kc��>vt��F�>�t�چ�	M�S�] ��@�1'����E���Cj�� 7��wjZ��ʟ޿Ѕ;9�Խ�˙�-x���[�+� ���M~���m�?I�J��ǰ����p��F0PҮ�y�>|��c�:M��,��a��1`4�0;[���QT%�X�
\V��YQ{�j��&�[<'ˁ���8&%�t�;������h"g`]�>V��fsZa9��<�b�M���WË3�42��R ��:�,�!d��VI�:�A��P*�pؔ�d���>���6-4ʩ0c43ئ�|�%��QP��T�_�p�
��-34�#�GqvuE�V��:��JR�]�4��`3�'C�,�9MX�ny$b[7�^ړ�l�`�
��4P eyVn�p� ��p[SW��(�