XlxV65EB    1aab     970Ȉ��7���l�E�3�0�r�AM/�~�� $G�G����!p��^��`Ǖ&.��~7�lsc��||��rq|E������=��P�z��:Q�5R����(�+� �����K�l�b"f]r�:v�.�ۜj!�;�\s�%�DV+� ��Q�e��7xޅ!�>an\?;W�ȕ�t;rZƚj��j-W�Y�|�Z��B��Ӣ��̬�m��|��k� ��� ���J?#�ҿu���NG�8�>8͗�"�	\��?Lwў��S
.��`p��.3,n7�Q�aH��P�*�����}�&HZO�~]4<	R��tm�cbO�8����w���?(��Tǩ0l���
�G2�Ԋ�X�haߖ ���U��i�CU)����V�TMP�N�K�0��h�I�G�G�㴫�m���N��z�����gV����Gb��וƗ
f���G��ޯ��7%�d�1��Qo�*J �7}��V�9�qqK0-���d@� �婻�B�J��^��Vu4$%���n�L���u�i)X���ܬ�A}�A�O��1��4@Z[���c=��M)��{zT��E�/9��wY�1�2�� F���nu���lq���q6�L`��vݚ�פ����@S�N_~�3�5f��h�_#�h�r����F_]n���ӭ���7P5Ko��o��	%�N�x�k�j')���mɏa�ku�� t�n��1�{�o��\l�<OI�����*��g?H�FY��偣��X���^�9�;\±(�$bƽ�����W���DC��{�����[�n���9h���2%��$�ޜ��{��k��I��r?(���)?	zY]�F�)?ӿ�"���O��!y���������F��Ы�����;~�	>Lw5H4����T�:���{Q̈`���,B�$�S��T1����X�h*�Syz�8��gs���8#*8�U�B�o<�?�x���ڄ/�diم뎰.Ŭ��A�]��߂w��B�a"r̍ 1��V�=������VE��(rv+u�����ON�n,(�7#Ȓ6����|�0� �VU�/����\i�ٓF��g�����'k`rh���p���7�!"�9��ϟ�s_�9����C�ܕ9������p@�!m��͵�V_�T���9�E�-�-��T���-��!}��P�T�W'��k���ώ�#)�`��|���S�/�"��ىn��!m&7{*�ġj�0E�V5N�Ax�����96[2��/s���/�Yf�������[`fm��ݫO�)��Ab�񰴈�Rm8W�b�r)ɳc��2��a�TŁ�$�m|E^>~�d��D��z��۠�ϣs�(�������`p�|c3�%s�>6�N�4$���b��O&�0�4u �.pq2]���j�5�(�a����Pf�d(:�r_���b�|n���R4�zt�����HnL��-�О�cB���_ z9�}��"�L}.4�U,�;��j�椐�}��@�[�nw=��!��/N.��_��A��v�R���w�Gc�⢁H�[(��V)���]���09�I!R,��*,�/\�Ma���Wp5'���9\�X�B�\!�� ��C�#�L���;m`h�:J`�t��Ӄ3�<λ�BI����RT(��(&
^��ٔtt��%���I�5�bJ6e`>f6�4�$��s	QG�d[O�u[�D�m���;��5u�ζ;�c���!�Z��P���I�~�]>���S���ڿ�}�]�H�2� M�X��i�__��6���c�ݏZH�v*q)�S���N������Ǆ�b�:S����*���"�@ٲq]�Κ��1fe9-c	j伏1�mgtu9Y�CFKh����Y�[y7��N�3�_�`�����6�%M�e��M���k3K���;5�,N,$�	�V�#�D��r��|Pu��\��柘���B_?��3_ ����>�L��//�A	��y^+@�;�qMq��a.#3���r:V�4=H<�&^��J�����\g0��{����ȳ-D	8�S�U��ST� �o�x-л���^�esq9G|Y�������vǑJt�,��4`wyZ"������
�186�&3��6�Ӛ��kk��p��� o��d�2���ne���*�DU���9�X���0޾����g�V(F��綎X�[�Nq=p��������J�j��m�t�s��N^ѱl��8Y��8K�����~S^×M~.Hl#�
�?x��A��ú�ְ��$�|�&��31d�0n��4j^-�Z�� ���A�*w�������R���f_/��P�z����cg�E�j���I:�7�.s�.�μ��M��Γ9Ah+#�*