XlxV65EB    8095    1780��yG$��I�;N��2���q4?ru�l����^�Pq��B��2��%,��{���o��S.�.�5QOPy�BhO��jh3}d�;�@ ׍a��hLS��u���]��bW�IN��끐�$,V,]�����c<��)���Q`�i�;�T�]<g��/�����CK­��w8�j�.k�Ъ��?Zv[�td꣡p��,^P��ʢX�xh+!���5>t����/��'��$��p��G[��C,�cX� �t+�;��Y�����z��j=�{GuU�.�%����798�5�위3I=�T��@@�K���M�cJ�S��LЕ)��A�p=�u^�L�/׻�8�;�'�I�����!��~r��0ʝR�P�9��2��(�����Z�_���q��X{��xZ��I��y����v߲|�s�N�S`)�F�#�![����� t3�k��B��v/��	e�.��,�cZƂJr~�9h���C�A24.�di��@��"�������N-{�[�=����Q��
��������Y($��FnK�N儀�U�������>��]�����վ8e��t�A6�1� Լ|:��Eh���Q<;5+iR�~ �涣�c0��R(҄##�we��OyR���m�\2���o^���!���ܶ)�ʋcR�'x��_A�9R��8��Q�~]77�H�~I��h
������s.M0�yB�n�6��~�pF�1#9$iD+�("xW3a[���M�pe���d�s��ߖ�_���w�M��B�c-��P+%�G�<|J����~�2K�3� C��!�7q�>t�V��s�m;23��&�3�>V��[<��U�°�BN7�C�YT��J���GK,�n�a�cH�0��S/D����p�?��y=��[�7�c�����W��!���
 I�6=S+ƶ���Ͼ�Z0� ���CQ`��&_��U�$��+�rY�t��*6ȃl���]�l)eQ>��D}n��\	�z�b��^�ૂ�2�Q�7���6�r@KN�z����l��3��^�7��<��ޡSm�A�M�_F�.�H�1}�`�`-�K��-���>����;:����D)�5��`b�S�_��("���:������&��������-�I���¹��� ��7݁7����҂Ci0:q���2;��A�p��:w$�W���[�`8+��g2??��3֤����_/,O�\G��^&�<R���5��f[��~���"������bͯ�`+�� ��3��J�!tV�g�1��{�!&麥��4�N��M�u����hi�[myφ��J�s�=�Ō�yu�Gba�0\ǋ�O���x����c�R�������ydܔ���
���M����F�U�KՖ�T�6w�
���W��9��~���g ��D7RZ���r�mY�&R(�OC�;�� ��6f�q�z���t���\�D(��u���o��x�=�|ԡU�, >ʸ������V�d(޳���CݕiSE*����]���x�����e�����uP���X:4~�Z"(Ne_��������a!���#LZ^��h�ižqs�vɮǆ�.E��
;+i�x"�G$�i�r?����bx��������!19��)�7�"} \�=���
gD����fL ����@�;��=�%��#��<��	1M��`j!��1%f&-#}(kΫ.��&ϩ{�:��r|���-�eh��G���"����Ih���K9$��*[?W�H��DI䕊��]4���g��\J����{>���
5q �p"���(tpO�Xk��i ��=���p�i-4<�a'��$Jo��ZJ���a�Q�#Z?h�{�iX�>t������Kg[�y���5�K3l���L9�{��o*��(p\V�Y¬��dP| s"[b����/r(8J�m��nT�B�������P�ß˹ih~��Q��Ј�R��M/�é�uc��wKЂ��5mV{΁Oϵ�9�ّd`;T'sTP�*^
�Z����I�)�/���QC-,����NU�oY����\�H
[a�m+G[���뮕�|t�S�Լ��*�~�)�?�/F r��o��E�G<�*�	J&�N�ZK��ֆ"3���K|q��'$N ���@S��M.�+ǿ�}�<�Ok�>Nݻ�t��Wp���AW�����dQ(�0�Lv&g�]ǽ�>F֧���F�=�����qz��:�9`��Z��+:����`Tr��-���δ�x&J+- �<Om�D'D's���׷V�%q���f2�(�J?@ؖ	|�#��l��ǁ�&+kB��"��o�r�������,��  4��h�WA{C+�rw�+:����\$[����Ƹ�ʘkA��U�/���I��W�F)��Bɰ�"��<7<HՌ|�d0=� +�A����~״�og5�ฯBn5��������b�z:���W�T�AD$��R�)gh��\�~��B��m�m��]<J0{�4RU3�(�\l����VG$�� �ȴ_�Om�H&��@�-�g�Uy���7ԙ�ma�c���d�X
BP���sg���E�Ƭ�6��:?�~UB;��A�?� 9���	L��&�t���$Һu����Sj�V�>T,��G�lФ�i}.ݹ[-��*��t�K>�kU�;����|Dk���B�>�	����Mt�}�!z�c���>ɫ�Z7p4<{��E �k�"�ES�y�>�����Z�^E2���*��G��;w�Ui��(b�P�r�������>�z\�U*���� �5<�.(�Z� ���8/��"�j`g��?Sg[TjKC������m����6��Pg�R��R�G��l��£=6O\���)5�}b�?h�����5j�k·|�f�x
aF��}~�������6���>��AZ�3L$6�(�x9�6i��G��Ƶ-�.5��*�Ew �vx���)H"fvV7�Gj�	٠�(0�;�Z�-s��<#�4ɦ���h͊�����LQ�z�B�<��K�` b�Jw39�H#�6�C�U�Rv^�C&D�p5������4f�ǰ��(�Ye��4�$�2�p��0������Ԡ[)I�o����/�s�w2�J���� �X�)Jv��tv�9���	��\��'������gt-��lm����]B/�T�6˯���/G��<��*�8tS~4�sL}��Z�U���,)o<�S؄9�cKJ���K�N�Q&�8�8bO�B�K��j�23�%o��u�0uQƿ��P����LOxQdyb)��7�b^��3HnDū��-3�g7_��״N1z�ȻW~��P�16��q�.��ԣَׄ�p��Af�=�JyX���r�S;�"f�}�B'��c���ڳb"�ܤ��W4��E�K�E�oE�����X>0@�'@lP���sF�^����PBT�L�ꕓl|W
[鵀ߤqBh�!o����2n"i�v}R���ں9�(]OX��"�Uַ��՜�j�'�$T�"h���W�S��_I3����㶽a����dS����Om �^�)-�}5�������'jfo�@נ9����]���9@A�h�!9<�|i���,o�M���=��ڗ��l<���R~I���3|1_n^k/!���?���]�Y�n�$�J���94̮��j�܆-�Բ�W��.��.����3���S�7]��DФe 7v��cA<#k%�?��lU��[Lb�M�[{-P�����'x�SM7D9�\�tC����<�Մ:���R3�^=��zt
��nS�w].��Z�����y��O��U��W`���Ȫ�F��b�Q����['�`�H�0��w���P`���`\��Q��G�)/h:��?���Q����$��K�q*�f#c�ʷ����\��4�;��ש�7^i�3���F�LA����e"5
(Y\��7�{�����b7-���T�+����֚�ڪO*��%hG.�`m.��v�uxҕB/��l(
�R@�H��P~���W�ԃOW������[��!Yő<D(މ��:�΅��;0M1ӆ1uN�c��߯�c����wb<ԭ,��Z\��ۜ�~��"J�/ZǛ�_>P���.�����{+��-��O�$V!�LD��e/	�����Z��M�(��7QK�=���#є8I�d���	ô�ίI�B;Ժ\���ǿ�ָ���� �t'/��nA@�D귃\�߷e���Qyko�p������W�n��`*���Q����ͪw�[�&��z�n+��+�����L�,}��~�A�ǜx��/U���D�ý��Љԓo���MT#_���v�����Ô�w T���eߍ��j�����µ
m�;�o���l}�.�K
���K[L�@  �l�U���5̖���|�I�_�p�)�?�����k#���x��нu�?�%\�%�7��f�5�*bO��h���!�<?+�hQ㊥�p��I'��8tU�^Y�m`��so��S
��$��;�:U�C1��;BJ�[�p��t� ��9�y��T�p�G�`O�F�x�yw�q�U}��V�����U��<�ÖS�I���㥀N� �D�I�*|���\t���d���Q.�� �Sܘ�Mn�$��mR����YJkd��0o�����_J�rEr���k�\����l���3H�~Q�	*e��.��EX)S�H��	b�-�����jbpD!�i�סt}�p!-Ц&6?_�27��ժ�T�^��bBRj"q4��Tt�;��D!�l����$K���t_�"(�'�#xo8��J������	��L�c�3�F/�5Xl���4E��]� ީ�/�S�WM�̄�0<�#ai�=�ac�?N�S1��6͸:t
ܽ!,�w��_VK�䀕�.��e�T�%r_]����j�ɠ�xEI6����(n�����^���{Zo��
�d�經���ã��,Ro�����>��1d��h��6��� ��SaTf�C��61C�vɄPV��]�d+�Hy:���(�`]-�p
���^N/��Zk�_r�xk�3	��
n;k�{��yTT{�V�[���.� yb=N�G8;�� �!7'�kF�j�b{��[�����+������)%!h)
�חg��2�RC"JK0[uT�m��.�Ȣ�O��'!c�ʜZJ,�7�k�R��Pt�|[0V+���B63�It0���
%\�}��2E^�N���m��c_�c����/]>�����|o�d
W?#�~kT�Mve�/{N�熢�ms�5�덭�c�W�5[^���iC��)�EU��;5�	�&����Q���4%ۃ�G��6�,���ܶ��&�:5�=G/�Fc4{��Os�-���,�͏&vpB���&���(/�i�.;{,/V�����-��8��5��oz�^>'l����g0���;�Rj�z��&dv��L�K�K|��[���у��QM�����6��l��1��������5���~AF�j��W<����ʕ*!$P��:����J1�z��TGܚ����]ᗬt��O��$�b�^�������s��6�<��a�3��)̀������8���̔�SF�<'�����n�#��᜾?f�Kp.ȧ�]Y�rU����Ղ��5�Ǚm�,����!�vf�1),A���Ȭ(�k�K7���PKO�[� җi��iY�Z�����QL`B��g`bw�X����U��;Y�,����DrH`�,?L��c�e��'���U�okϧ*�pA�7JL���Z��J*�� ���"M*�hO��p���Q��]|/��V,�	�*7�3,\I'BLW(�/��I�I��aC���>*�w�h���;%�B�w\!X~�+I���o`�v������
X���#�����,�O����<�2@���|�m�	3�|�