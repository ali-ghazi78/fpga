XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��n2�I����q5���*`x;�s����MV�a�H�ݎ��GI������x�(Vn�H��=���A���%|�!��L�r���(�e��6> �i��-F�MR��w��L�U�u!��U�~?��h&�L�5�ٚ>�J�w��Ã��T�8��������.K	�u��A�?"��u�3F��G�å�o��76��lab�*�ȩꔧD"If��N����>�Y5!B-���USv���ṄJjd�v�Ǘ��W5`��VFӪT���?��yDv�$�]��"����9��*-�,�����O��a�0
خ�7h^��?��V�8i��M}�����֮���As|�j�{����7FB��՗s���C�vG��=Hh���tҀ�G&�?Q������p�h�1`���_`���a�{m%�5�B�S%;�K���b<%�"�����/{��x>��k���`9&Н�� �p�	�����.^xa+�ѱf��7�˘ɟ��lB����*|��sޕ�T8;a��n�����I�N�]�<���'�m$ �������L1���R�$�V�������`��`S?%5٬���,/$@����8Ğf�L���z ��g�JHW�,J�/n���%2�E{O1ls����#�`{�p���\޴d��1�J���9�&U
O�
1���o�=7�n�9�Ѥ�~�Em_��]$�?,w>�30w�'Tٰ0@��A�l�l�R�'s�9ʌ6�	$��je�1�̣�Ǎ�XlxVHYEB    1aac     9708���V5��)$����СP�����|�Uv�p͒W5y�Z+q�Gg�GC3pA�V��s����)���+kBA(^�ܘZ藣a ��!���	�f���	Kzט1>�U��Ny��Tia��T,���d�$N�%�,ߵp����r���c.��?t99�f��v=-V�``9��6m����Mzv�������O4�tC?�yS.��1�X� ��<���W7���d�޵��� =���e�ߌ������IĢ,Vo�!ҋP�!W;P�������u{�U����*�?j�)6���T��C��$N��յ��;�Q��c��{��^k�aeBE�Ci�&�s�\nСܮƦG"6�z��Ŝ	����AA�6�V#��hQ�mӫ����x^ *�������g$<g[�Ϟ�i�}�a�[��#K(D%P��&L�S�h�+/�Y����.�|�]�'��D�sI�*�NӘ��N�_��F!=ȕ�5�0�H�}ʰ�y�[t`�~[9Y���tcԾ��G�`�~�wl���@��Dh��m��� ��oe@}E�Y>𸎝�D{��%'�q:��G?d7z������z���g�d��:��}O&a�!�;E��T�c�$<�z4?�tڲ��֡�>�$!��'�Ͳg��9��Zi���Ċ��"LM}{�_ZD�FpI�)#׳���$n2��XOD>�(G:��,ެ?�֦i��x��*]��X�R�a~f��^.2}`�1������r'��@/_+��gҬJ�k/
_":��Ϩ�)��t�PQ#�D!��z>���lg�.��VK ���*��{�h�A&�e1{BMb�W�0�,x4R8��|��#NWH��1��D�]X/��]�v���R����W�.œ_cO�-��&s).졾Py�@�c'�q:�����_�ۜ~j��sa7Q��H��%�����iϽ���:�p��!m��9K�]�Y�.x�r��}�1��r�eC�7,-�x<�"�T�,��8�r�j�;Hj�/�W��Ah߆��~���<�Ƕ7�S�濇�� {����$!+��H���t�.~O��-�6�����z�$�g�)�:p��ãuX�A�Ym��*qƨ�b��� �^�iR�Q���	�H���mKȨ��(j%� UI\t�E���H'�2r�!A�f��V�E|+{�j~f3��>\�Ƨ&�G@�_�z��BR���`GŃ���4�y6���5���](&���~�<�.
���PDN����'QJiQ�W��u$�D"��Kܐ��DkD�}u��"��Ծ3J�:�Z)vf�J�Ú�/K��?ڵ׸n,Gg&���3o�_�1ߑRcV#��7T5�yi���\K4�iN&|��.�S��}��
�g��0�<�sa8!rzQ��S̿8`o���z��"����'�A���2V0�{+�#
_����Qh��4�b��{\m���ρ��La*���>�S��l��%�5�B�c1��[�YѼ�T�9����s;��Fֶ���+��tq�1><݄9I
q(`F��.�٭���hV��z�G��d�9�ʸ����1�N�uҩ`p7����5�78��ïE��2I����a��G��(#��_���d�n����E�mˉ��U
`�\:_{���)cŴ�\��.��
�B���e�4<�9fx^٩�l��B��*5��ﵝwv��!ױ8[-r�d�+�4V�����T��0-�ÄÂ� ��_�B������!�ː���t���<���:Q7������m�#S:��A4dU��z�(��iq�;`;�8�����n�O�@9Oll�"�^L��Z��.�:�qO�T&�D{U��V^�����d1�9�ۃ��Eخ�ˢr:X�X��or�-��L/�l�ҧG3[R\0dB.}�Ҩr�]�	?��u�"���1������N~P+�=D)A�#�9���)q�����j���V'�/��%�?�IH�~M�ժ����o&J��"�5�4=}�潌���%���8�T�`����9�h��mdz.�
u�,�U�V�R�g��5����|�60�O�e�Z顀��m�o
Y��A�g�e6�<l���4�����|��\X�nջW3�#^����B�1Z��C�g�.�����mLT���:�C�f��,�2��Cv�o��M�IU��L������m~��8虋U*��N��͒��,�;wS����@�7>�ݜX*�8m�aL(mᜂN���Tr�t
��`�Ď{8A�c�D��|
Fu�bF �n2B���P�m�I@��#�}����Sy��=���V�7�4{��U	Y�a9���i^�+lxb��������2��0V��o0��'�=�<˻�{<��]8��-a	���^�캔.�C