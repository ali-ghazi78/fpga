XlxV65EB    2a38     a20��Y�
$e�$����V
<��ӿ����C2rZ~@�bt�u�1����US���8D��`����ږkx��17>��oT����2�lUÃ�\
пe�IȬ��.G��ߏhx|>�s[1��͔�F���b�_���»�y�.�nˢ�s�tѮYEAQ�$5*4֢R�wmh]�8Z�]F'��U�g8�|�](��@!���[{^����A�q�1�1�7��08�l�:�T���	���@�5s�����m�������q8��I�TT_��Nm�'x��L�!v7N��f�*�r m#P���W;-���Y��.k�Y� �>>s_����j��cs5��~����Ki���sⲆM�=Qv�#����X�(C��p�U����(X�ޏ�a�v�׫�f���	Iy���*��\��cȵ��m}_��S�(:_miBd����W������$%����-V��)4�h��HO<p]�i��VP|ڌ�Ce���Y6���D�3�+rF'[��<���i���-���t�3�鑬��@�<��Q���5{e�@����zC�Qb��&���6��>r�ߴ��չ���U�xd�s;8@��͚�y� "��8K|~pD��%�#��14]0�JE�-��"*%y�g�G�R!��Je�����1�{d�Ѵ1�I Ay�I)W_�%`OI�i>��]����_��=�*�����o������2��$�]^x�9�������d�����%����L�,�v�����	�g����,5TQӷ�9�CA���W�:��ݐ�I��^�&����*���R��<.�V!S��J\&����^v�1�D�W�=�%��zR4[w3w`�p4;� ��{k����{��U3LJp�[��We�8de*�6�����J� E�i������7.aQ�_N"'n������tK�s�7a���������+]svY�B=�^���nc2�H)/��4��@;.S�����$Ï��r$	d��q'h%k������t��X�Tn�w��.T�Y�2ßWҌ�?[�3�]�(Р� ��ku�kd,IV���\���3X���|:J����lh8�bۋ��QvU5��Y+6"���bp}`���ذ��/� �Z�4C�ԭ=�-�P
�˷*?����Mw��

3˅Q�sx�*��:��B������f�|�Ǚ�N��!�7��
ooȻQ~���|��� u�FNV�H�_���
���n��k]fq�Ěw�C���J����*��Ѳl����Y65�Q�P-lC:��R��U��o2ݵ�!/��?_�� 3�$QF��᫳rrL���܌����v"�eb��+{#�<r��7�lΚp2�t�� ����G��h�O��)�J����d�ԷbT���Ln��[P�G&n���	O,)|f%H��YߊWr��o��;��7B���� H2*���9����H2G�!��nl_Zճ|����Q��0�����e|�!��{y��h���eL>/J�Q�����T�����w�8�Ҫ�R܄��|NC�lX�K'��6�D��Si�\ŅtH��k0�,Wn�A��q�p�X���e��no��<�C2ʁ(3��և�n�����e��)��B�;<��X�'����a�\-+Q��J}�/�X^�w�U�R�"�ͭ:"o����(��U�tv�W��R1y��(xR#�Dx]�(����o�B�owB�� U�C��^�����R(Y��|/G���J]��5l�@}o����&�� a�Y��-��Dmý8�Od�à5���>�/E�[Zj�����z�$��m4�zQ���C�Ơ��@��j�7u�mr;_����b��� �k�i�Eq"��s�Q�؆�[�Ԋ05�'q[�Vޅ͖P6n��%��>��m� `e>~R��J��ׄL�м��ܚ��N��6nш���=BB�^�V�j���Kx�Fc�\�b�xTWE��0:x`������R��s$�KH�j�sPֿ�#����d��+`�ٰ�[[`�:R��w��SnX�B�E�ki%S-���]3?~��e��o�z-��B�!��=
�E�;�q��ރ.ٜ�=_~E�A�p�]\ě�+�f�߻�MCQ�m��)/l�kwm`�5����7%�f�Z���V����(
)+jL	K���E:��%�����m���b0�aĕ�<�N��U�k�nnB��(�����Vn<���M��En��'��l��;��[���k���L����ʦ�pm�kվ�{<�0��������>"B��O��~��3�6gf���殍{�)������缐���f%��\�טy�/��F]���5o֞�r�{��;l�ҋ���� �:�e�Q5��.@2=U���G�$cB��I�C�Dy;��SV�KU��m&C5b�db(�)r��JBt�8���14	9}::�m̹��d0q���A� 5����-8�����t�<5�C� l���s(è~�_g�% oG0UN���P{�7�������(���w��m��{�s-f3���\�����