XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��\|Zyb�HZ�%��`p��t��T�Z,���n%F�U�xac��D��+��p|��j뇿�Z`0��� ZXO�GM��e�)ԕ�ɓ�+�鶐�U�	e�Y`wڟ�:Υ-K�BhY���j������e�R4�JMDS^��*�n#L	�hUA� ^'+'1$��.Of(�mkr�Vz�W������<�"�"���_`��a~|�H�/yu�#~���E�&|p���6��%O�o�ݸ�X?�&ʥ�����\��0�#�d�5U:�?�y���j������� ���������5N�D��/bs���������Fm�:N;��T������R�W�	�k(�+{��X"�@���_��9�Z����[���^���貀Z�+�H�q��e��fR�ы�Wȅj�L`��a�O�u�
^�2�O�a���'	�Vw�a�?���J��r4g�gzz �ቋ��(�^��L$^�{�#����}%^���h��U?����;:����#W�`v�~nrc����Z��w��~���D �s�"�4��/�VO�sm�(q&�*��a��ca���ăXilʇ���R�F��^�//8�v�1ZErXۘZ�����Q�K%F2��I�4�>�݌�aw�;�lIKv����|Z�d���(#��ИJ�"�m���v:*B��eE�a�6I�˝�޾�˲#�CC�Cj>�Z��GI��!2�/#�@�Gz����_XB\	�F����.�d�~����(0��g����ur6$�@�XlxVHYEB    528a    11c0
�c}s"� �D����V�����ǟ�0�
LUU�飻rX��r�ݵ�[�W[Az6�T�utɲ[����o�3�7r�~�l<3�*w�U���
F���C��w8�^��9��U���nZ�G���%&��_+�tˌ6�z�h"x���:��Ĳ�J���n�qȲ��Hh~$RdW�S�.[�x-�_�N��\S �9��׳�C��]��y0~�+���w6��,�ډ�˻�3a�Zժ$�
dq��I�����@J�H׍������('�a#W6<\�v�7��፡,�����Cq`�@Y���3ʦ�ژ���89*$�����J[8�r��R� �\�cM�3�,�?�r�7,D��UT���Gx"��~�(@9��"''B�X�����B��Vkӭ�֟C��U+��!�q�͘N*�W�%/	,$BN ?�)�L�J<i�\]��$ݲ�mU/ط���y�+J=l2�]G��eS�Z�3 "v���R���t�3����x(8�ӿ���0I�'�k�Ws�2���M����0�`��k�r��ZV�ok�YE-�L4����T�Ά����S��Qe.��㜾ѭ�;$A�1� 0 ���?"���k��d�!�k3��A��H�g�xx���i \t�X��v��buf�1���a
��B�R������䅾,��5'�c�n?�ܷ�����7<�i�ݐy�
gO�vB�,w��@b��X#'Nr8�3T���AOP��Y��Fzi����Y��-��s�W�}��nĮ�,�_����'C�>B h�:��K	�]gK��]�;BΠP+��'��{۱E@�n�MU�
�C�Ir�SM���w���|IMV���
QC�9�_\�Qρ��@ؽ��u��2��ŧ���Aq� �o$��3����e��tl���e\?ɕ2�P�	'ڹ��Z�<Ő��<;�X��>3B��.!
�8I�0a��W���X�ٯ�wClDA��L��<,�0�����XK����Y���<��j%x9���L"{�F�.Mԑ��qQ}�Vt��v���>����%ċᓹQ�Jn�oo0��Tۓ"��ոDl���&���IgB�p���̘��`x��]y'>P�n9���=Gz?d�V��5#׶��Y��s���z�zhZU3'ir��Ͱ�}�p��l�.,r�b0<սO�8��F�� �K�U��w���Gm8hXg(��ճ�6"ʬ����W�cT�/���?�mн�1`�̲����V~���G�b:EeR��}8fv�`_ωW;��c�q��Kzzđ3V�	7/�M�2%������Y7��iZ�����4��{?�j����8�����X�u�	3QLA!�2��nCz��5B����$`�H�+;�=*|�[x_%	�=��1�c2�f	�L����A�`���6�L��狫����n|'�vx��NVg='��u ]�Ke�?�K���ՓxR����GbA��=N��	�]XW�L�p�M;I�.������bü���?�4D!.t�w{m��R��,U��s�^��#��\ݽ{�ǩS8��'�jձ�d�k��&̈́69̟������?�����������q`,7�gN��0t���JGM ��+���������)�g@�?�_¿@��Yħ��� �0M�������RT&��N��*�lE0�h��
���}�2�a|TZO�J��4O��p"f�R�6'9������O�L�#��������[Q���a2�&�^��Sؕ�u��a67y�	�yCh�6-(c2o�me�״M0���k1~b��;W�9�E:<��^c�H�ɵ�"��.�:d`���Mjt���[�����P�-�x����R7��B%K���(o2\/�3�����s=xfO�s���mE}	v	�&�`��'�<����	>�k�U�8O�~��������mp8HXf^����G��J�ot���ӂ#c�U�3�������1��M�h���C�eٛ�8.)O��b�*&��Ylٙ�4�4/Ѕ�p�
/��Ө�g�f���I9&fD��F�v��+�qD��%�=��=�ʦ��8�`�bT�%���h~Y�����N'k	a�>���RŒ�3`��J��19R�@��m:I%�E��5Cfi`����|f��"+;8}I�('T6��%����6AS�G/(�ϖ�B�I�4��agz⇸�PU�@�"��.���������a���hA�7�����+�8�L�����M3�'/�{�K�O�,C5~-�i�O�Y��SQ>���r$&�'�L�6宓������3�_��&�I���4[�Q�$�ІFgPo�]��:R��7�~L� IJ���ѧ�h�L���@�H��Y
*{���ߛѣK;�\Wס~�:
�F�!v�5�ŧ�N������s��8����I�5l�Ӏg��)�5���v3�����[^t�.�ۤ�B@_4�D�Տ�K"�O�P�gk$ER�1��X���aM*of,�mH]�g6�oP���,G���q���.�8���d+(��OΪ�������
R�{/\,)���&��:�3-xe�9��CG�K��[`? �D'��YE��tmP�b�E���(��o��yb�CI���%(�mJ�%"|چ����[�=mҿ�K�p@��h���{L3���W�]�L@�o����{薬�k%���b�F��9.�	��l�.��LD�Y{v�O�$�3\Ҡ��t�� cŬʐ�vsq:����2%�
7}Ľ���ON|����=�����գ~p��(Е�=U���V"����Z���o�ZaZ������g2��6�Ԍ�bK�0�ج{�j���G�C��2�� ����1�j.�i�!�<k��;�cjoי�ue�N�Y��6�-�h�=J|�`�����Nd͉�t�9��1ū%�ִMx}6E�5�P3Bp���x*���1��ԅ�nF3b��_�ɸ��A:��p�}rHX��nX�(ͩV��gB/˾EdW~7�l��"Lu����P�	r�V��)M0����d|{E�hq����!n�3!������OE��Ż�d���%CD���P�c��$��$Y��6�G�W�ntL9�����ye�`
-O9nvJ'����7o�g�a�W��ꀜ�t����nXXaT�e��(�f��Z����8K&v}=g	���yǯ���-gt��>�G�`r�o�GQUF��*F�--o�,���*�d�~����=�{��͜F]��*�$����S1 �k��"Џ�������	k���%h�� 4�Ę���%���v��F2�����?��W����t��J���;�5b�)_ۅp��semݼ�T�H�Tkk�$��G�ru��.�wJ���G�23�i�ZJJ�oN��ty����-1�U�"��NnPI\`|���g�!�� �f��uԻ���pw�1s�� x�ʌW hz�����2��:n��H"����_�UM���ۉ.���ȁoڥ�3�j��G3~.Y�I9E�pζ���rXǡ�6�E	��3��M@���#�:�:��1?�@���N)�Þ�dw1SrK������7!6��8U[[��'�{먱A��c�̒�F[��v*l��	a����'�_���h��2�hG}}Zu���2�q*!�֘-k�J^�?�%�2�'������[s'6t��c^!�������*�Ιg��j��ǳ�hRb#��!*d��'��U�*���:,�t텖��$�߅��-�9i{I\u7)}uN*/+El�k.�O�l¥>��skF�>(�F�u��~�S ���4E���b*�9.m�ʓ��
P��91[6�$$�(�0��D�:�D�T����!�C������D�4n�ޓlQ�I�732k��
jt�[�����?�2�)�D��'9@��d����s�ۑ�m�RS��Dk �Wؽ���z�`�A�:#*�k^���'>����爱�0�/��n7$��1P���뛀v�z����c�$�?�%�s;[wF`�ϙ%:����2[)������f<��G��c+T�d}���P�;�՞��i	�1i�;�5LW8�	�s\�L#�I��q��H���5����/�B\Tl���J3O�b�����*���2Ad�K�-����6�;a g;4�uonM��\�¿i<-�}y��Rc��t�
ơ/�B���� ���p�L{H���(�G{G�����/��fS��;����wZ#a^+�>�^��� CvK��:�*�<����7�-���P�֚�x
�o��z(���p�DdS(J@�Fl�<V�����"�`SQjR|od�h���S�]���2' ¥�:�~�� �r#D����e>�^�"0ʆ�:;�l
Ы�T�Z�\Ydj8XJ���nۻ��)�~6���&9���xѰou]�9,���T��x���V�\C���Z�S�E��