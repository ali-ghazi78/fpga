XlxV65EB    dae7    12f08M�_'�mj��c|����n�+c|9�zJ�Z�,'���HX���p�n�cϵ�N�&��>!e�*j�Mܽ�1+���պ�v~�T�>yh�tl��c�F���$�8Q��� ���f�c����E�Z�$I�2������A�3�cr|\��،�5Wc�� V����K#��Ŧ�ңG����mE)\�C5�P5�9Y�.���Y���h�p��tUK-PM;���vY��0�;!m�� ����^Z�T����Ϫ���*�l�)��2L�gXjf~���5B�r��`���̴�۞��/���:�&�xU��/3S&�O��͢�&���Z uAL�,ֈ"�
�����e��	L�"?ƾ���*�S	1CV^R��MXa]�&�U�ʏZ��OD	�>xI@kP���.�ݡ6�ȗ�9���R�|�䤂�����%��
����@��C/��Q._<�ש��W4�C�)�F�zR��ŵ�pH�/��G��E>��+�d:x3E������~���+�껹���;��N�R�x=ߛt�k׿XCy��s2͹XP>�P���4���Ĩ�+��*0���EgTU`Ļ���,QK&Cʁw#��-m	k���_
��`g���A;��b[�w���
)
xg�K�,n%v��� E�i�U�bh֎���簕l�<B��:��óL+t�| g��q��C�5I  En@HR��7�Uv�q��ɟb�rtJFA�t@m
}�e���)%��c���4|į5n˺��|K%@��2ƦH�o(Ҏf�D�8ï�	(�a�A*��V|�N����g�����*�1��x������H�ڡB�>����e��R�r&��oO�Y{�� p����L�1/L`ֱ���������%�������+�j���>�O�f�)iw=� K��a�oN�[9d�[�
�c(��ɵ,4�js�J�GLZ�s��7��N,�δ�+�����zRV�kF��\)Q��i(�ƿR>]T$c���7��β��"��"!��tpa0������l�T��:�Y���4+ah����r������ʎ�c�L�û�R�d'�1�T���p92��
�l{�V��N��ǥ|C^k����A�!J�-�	����[��B��1
�:-�7���Cݐ��s�0��o*^� ����4��b�Y�k��pt��Z";g|�-_�m��GAz؏t[�ɂ'���1�8,����0���Kn���[m���qK��͘[�����$�ś��7�P�t����$��f��a�*��emfR���S&�Q_il��U,�	>�v�͵��	�&�䚹3�wJ�u�G' I�J���� ��1��}XxVY/���=��(XPG�x���X�7�<�Ba�y��^O�d@�T�qxP�w��@�B)��B�S���~�d���_�i�ofb�L���;�I�<w�Z����o%0�/+:�ؿ&��(�T�&���y$�.���U�r��I����3�킮 ���s��lq���`�U��P+]�+Q��/�}���}u�W�ڏ]ǣ�dL{U.�T�L�o�H����z
F���y������f�� Њ1�⡑5I`�x*�E���1t��"�Ĺ>U�:@�n��=p{��>O�/bz�6����8}�w���� �qG���I�
r��F�b��1�R؈Sx�7�i*�H��	�DnqH�j�����A���^g��F����zǶA�j}�P 4��6��`�P�A ���  F٨
\Y�,s�0��"�|��򛿂!�v���k�z�\�]�!�`�{ʩ�S�C�!���>y{�����遃p��0��]�99�[�Bљ���=DE��y���pQ�͙�GuzǶ�-EOZޒN쁵�2�`�!�λ�y�'"��i!�>��Y�D#�AX�b{z=�_9g;���A�����SX+���&N�a��6�n�C]=�ӓy6-��\b���݈5�?���͋��rb���략�WR��#�������=V��X�B$m_ź\^*M�|H����˼�z\s�r�_1ވ�29 s�b�yÀ��Bt�R�����qI��9񄥊�/��!�@*�u���wu�,!<fZ
$�"�$2S3�����r^��_j�f������u�%�L��s�TWs��?v���*��Y�+5�˲vT\[GI�C�pL�X(���8�N� �:ŕ,T���ڶ����9UR0�����k��4���X��jziצ�]�G�k�x�����(o�^_�ΨC��.nV�\�`�[���o�n�ر�F[-�zǚ�w$�+�4B>��sVz.�(�a�~�W׈I��qV�BIK�S�fV��S	�C��8[\�m����K��8@�BYױ�s�7q>�No7������]/�2t�	�߶A�t��hx�_����@�uI��Bb�n�[��xQm_���P�6&�1)/\`0�
c�[U�y}JO&<ps�pV�M6��)L�> �wQT��I���1��lI~Ѳ׈"��L�C�ul�2jX��LH�'AAY �Ulo�5�Wp����͇G83��>r18ß6��I���s�L�wQ��6P��꾗� �v�(��Y]��&Ъ�n�s��4P/�!��6��H�:1�M����.��h�bs��������]�ܒ���>A�3����i+AJ�#�:V�o�T�VɸyC��u���224��ky��P&�����{,5|���q�3�&�7`@'�K���dX<�$�����ڬ"�`V�X�F3X��!4�V�U�! xSD�ǽ��q*N���Iʋ��E��ZQ}��	�E��N�K{��bYe�9pu5�`�'���*��(	�G��k��M�IѦ	�3.�1N)�� U��;Y#Wl~�j��,�P�ƖLm	7�p�����5���S�+����6��y�W�h j�F7�|��A���I��z�oyĻ.�Ac�c.�ḏ���}5�|�f}"����?���`��ެ��0�ďkC9��}�ts��L�	�I��Pu��)K�����g�"�^G���ĺ�J���L���"��(u����.Hr�#�-����c�<��F��ۡ�`�+%�|Ck�f:OAd#Ņ��4��@ݐ픯�Y�_v�HV���6kS�Yw��ikp��&�/��v�EC�lȬ�>~o�K�J��H�Ds�H�a*����[�^�K���4���V��{�4tC�F7 	�o�/PI�r�%����@Z��QKlػѓ�u��A��ʕ6��(��PG�dA��l�γ�!�i~�6���Zx�s�
��}#�Կ��T�'U,��h��\��(��dR�{uKc�7� ���W`(�3
�3^��/l[���'H���v�NT�ɖ�����̽ʱ���ؚ��>��)��XJe�#y���s�xK��Z}DEd���Vk�3�a��hn�i�ew&N�v���Kc\��s�L�?�� �8е�=�$_�+EH�B( �Uc֔
�a��o������ѤCz��k�zd�c�wt7e\"a���D0cXhN�R���d������\`!��2v\�F&�%��Ⱥd�tP6��i.L!���N�W90,y�����R�c������ss�c�F�9�5���
���f������[��m�!a�R�s#��: {�����S��ƥ�h��j����µs bP'�������@��W��L��q�� �F|w\<Oa���糱^���7��v
b[**a����>��!���IV���6����s-���n(������2�W�d��ύg9�p��^c��6r�b����\�� �!�R�����kUj� �+oT���#0���$R��w�@ha�O�i�����E��&	C$X%��ǡ���es,�_��|}�GU ܮ-�:��5,�{
�\W�3cd��7'� 7V-1\_e�t���k4�B����N��i�����?8�Z���R�9Ms�*�U�恘������*h��R�B39��L*�~Ɵ2�j� ﮗ�y3{�}d����V�p{�<� }�w=Ӵ�N���������|���Ϡ�A��#�%\I���P���v����
i�
��w���g���Q/!���3�>N*���H�P��s�75qkA_� |v�ۇڬWM�t����N�|����"���o%�(��vEu��!��]��]f����$��j�#���N��t��V�SJ�����괱�dA�H7WU>L�3�ssC���m"�𕲕���Y��/�!���͔�᪡�m�\�, �G��m�&��߈ak[DP� 0���Je�Ls��ܤ?g0�~Gp�.�y��2f�b��:�[�2��6E�5"�j$G�S�vX1�j��F�gu�@�Os��	%����@?��%���A�:�#�qJ�������9��v�o�K� Q���!�m���5\�=e^3�;S7��G�T nt�W�1@�x6̗��C�D����?���+`|��{*��k�C0M�7%��7x+.�8�V���C��`=�ʃ�u(uQ��G��jTP�:�ԩ�vA0H���1�37Y��Y���}�dCL�GE#��qe$z���U֊��L����̎@w"<���f�%�unv+'yd���/ߢ�SZ���.��tg�������厬3����HU��u���0������S� �H��%ɲj�v#����0o��,}�@P�'��z��s�@ת��� ���s_�wh�����.qD�a�;<�2R����0���