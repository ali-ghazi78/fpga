XlxV65EB    136c     800�e[{_f��	,T������y�#�ƣϘU�QZ�B�R����d0�h"9	�@�5���ͻj�]�J���Y�?�eEKV��иT_�x��mI+wGՔ�i�8��~y�[�d\��d�����-�7��!���F��Z�S�(<���� ț��XV�Pv�/�WR���LYKMch.��ϋ�<��W/�,m�iDX��ѿi��6�ҍX{��-�t�]e�z��or7!��$i���qW���"���0טNeq�TK��x�8R*:#V�}��UG}�v��A�Щ�#F#�����|�`&�	�(���p�3�WDk�LF�>���؍��O��_l
qV<)�G�"�@nq�h?�uϬj������=��C�	|Vk��LX��
SAw͍�Rf$%�!$�:1�۫*�v2+��x}�|�����F5ˢ�ԚwuS�Ji�ϧݒ������Z��-��n2V���v�6�����$#����`rr\��zO�ᨉ�L�{�=�ή�	�h� Z�	�R����P���"X���n�V�ڦ�������[�� R�Z�'�$׳Hee���{:���!�˳=�]^kR��B� x�k�<�8�'L̜cq�MW��m�gh�!ɺ)&B�k'I쀛?|]j+��E)�v��i���qD#f"�����d[�a��U=�Ӹu��u�w�z��4��lM���$�$0��������f��(�Y�Y�]@hԑT��HkN�����6��M몿�����)�5A�X�~3 ���	�F�r.�U�_$�[u�����+6$D��I��'��z�h�E��Nd��[+�n�j��:��Oy�J
�X���Z*p���\��Ed�m��r^����:�9���)����Ҿʹ�;��kCN�T^��Ji.C(l��k7��N���<��xj�����KR�%?���赧��f�e*���?�ǐ�
o+�x."�z�]T����?3"�?���o���W�l�.G��R<f��m��wK�>W��1^;���`G�P��N�1���s��q�"\6�7�圶���$�CF�ki�����}�k�����t��Uʠn���eؾW���0.}��!$�ʥ:#��fꄷ��!�"�-V�E���,�����}a��d�V��5k� a�t#�DNs3�I0[J�@��v�k#�ܖ�=p�GDtL�R6� ����V�g��m�7��������V.�0V�I�� T�~�%��-L
u�v���n�)f^P�pt��-,V�p��m"�*Q��Y�㰻wr�ŉS��%M�|/e�U�̇39n��~Ҝ�E�F���õƵ9�Ԑ�%G��Af�����k`�f-��4b�'+L���(�瘁�M�����C��ɒt�Z_��{�P�M��γ��{O�Ez�g��&�y��+����|���Ꮆfhx����d���+�ɃK#V��N�K�M[	��wW�o+���y�*r>=��d����V��Q�ΙZ݅�F1�kbõrQ	zF����誅 �`��
�y�)��7)s��j΃?�W�ΑO��g�^�Ŷ�u+��r�
�fO�K�d(S��2_��DVg�플V�����"��rP�6ND�f|���td���u܎/�B)`�Sd��������o��M�x���v��g����S[�}�80�}��>�����N~�5��{�ٰ܀`E$�cA���
zy�h��b5٧j'*�I�+�i��}Z_�1ә�H���rq<�
��	x�>��EL���v����j��Ry�V�V��<����a7XC���сt^�R���e8� �?N'�D�֥� ��oӻ"B2WG�uV�m[S)L}�a��:��"ԁl+[3�p��xגB2ˋ?�,_p�Ø�������0i��2:����P���L�1r⃣�K��U�x��ϟ����1�x��GKo˹�̯��4��#���X�� Q�KT�Xu)�*^����ش��\³��r �hf�U��J:+f�E+I�f8�\�J�V���W�