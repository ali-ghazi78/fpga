XlxV65EB    1a28     960��V��3th~���^�7��g�ۼ�+;��e^}���t����O�=�s)_y��隿kOR�����"��E,�m���C�+�S�ϣOy�1s|����u�zn@�������� �%N�4,�	�K����2�F����� ijl4�Y+PiɎ�\�O�t�Ǯ�o���>g�C��`#����!�H��NZlr�v����["?���tW;�#oL���&7����0il�<�$�fŚ��u��ܐ"�{ 3���У�}�g�|��P�l��N�Qa���Cm.1a!J���.�țZmI��������p�dAd�}Q_�����h���1ت�\ڂa����
m�9鐛�D� �ɋ�r?�N�#G:�x�.�ϴ�ҫn��{�ʭ	�6�e`�����f ����6ώ�}��_���i�H�c ��]�cMq{x�}��6^\pUZ����� ��y�u��ǝ#k��-��T�4�PhjFV�g2��W1b	|�D�l��w�X�/U'24�BKU
��ms'�86KB����>:��v:�FKF)3�t����Q^�%�T|��8f�!��T��v�~�%Z��Ո!����A0fV�~�ga�p���nrܞx��"��I�;��G��8~�����Rvs�-�a�*��BH�T���Q3dU�,�26�� y?����_�=������dP+�_�x�]�q�5��rz����RKts ��)�	:`$�6��&lL6��p��G��� k���$��dߌ�k(+�R-�w�*��dw=c͉QZ���#o:����ĩ��A��c�b�l�H�J�l"�(Q�%�_�Z�C�����`��	�.�j�^�ĚJ�dm0^�O���f?�*D�[���YF{�!B�����H�6�B�����	J5���/��`�Q�e��uƋ��ck0��@2�I3�4�r�B�^��@�l��ǝ>+	vBbx����)��Y�v%@Q�}1���R#(�å�f�Q>4�ި�q�0�U9�����xk�,��O�.�θ:�G���pĬ|���ʒH����)�����%�b�?�́���g��a�sH��2�9��y��A�d\���T�C��t�:QeS�ܯ~�c�@x�0XI	�@���$�J�����G�s\�1�� ���i��'��,_��_�y�$����m�)�@˟"b�o����fh�pV=o�`Dr�s'�����h+�a"�Y��a�� ,���v�غ)��!rOxO��W��d��㩺�i���	�vO�vʁb���F�C�?L�t@���{��,xG�LN?���g6y��[S����"
�����0U�Zǌ#�����CNn���&QU�m\����ah�H�f<!�\N���KV�x��{�<������hN�}k�J�$�<�h:r2^���M�GZ{ݶB��Yն�h��asٛ�c@�2W����;f.O��SP/����u�d
�[����y;�ՙ����ْle���X�5���H�����_�Y<�E�1�h��s:���v��}�=�d!V��ۨW��l��=�@����"6]���H &�F3Ǜ��./;NJ+Vx�a��J�?,�_�U&�	LP�yl>��c��0�l
���8}7q�^ȿ��J0�E��u�M��c= ߫;1�Ѐ�A� ���b���DAj$_�t�r6g'm��!�T�(כ�*
	�t�z����+O?���
��8t\���O8�W�H��=�;�p1����ǌ�zf
6�^3����P�j���<iB[���d���	\Pac�$��砏��}�ȃ��S�ez)'"΂H~V�/F��1��OY�?�0:D\�ó�o��E������S�ٌ��֪���^e�xz�J?����HmÏ�|�k�kE�G:[<A��͸K��l�-�cA끥s��:��� �cZ��̩jM��cJU��?̀@z��\#{�(P�!	~���M�W*��F��:;��x�>�.��l�َ��ki�.����sղ�f�3�
�n���N:�G��d��Z�����sS��[���aL���fY���s�5��w~)娺�$�`Y�K��q6����2.�ǟ��wX�5��F�q��P���Wc�eiYy�v9T��#��:�ܖ�>���wCN���e\�S%1�4f�$�p&��rьĠ����8���Z+�	Ru�6 .6]��"]�r�������������;2�Z�ތ/n�ȼL�ͺ.gb��Q�+x`�5���9�V�W旒��3�W��4'����׼���T�
\w��``�I	�gE��Or�}E�hR���(O�� �%��-�`k��]A�U-�(���:�\�A��K�KΟ�f	�ɠtb�O