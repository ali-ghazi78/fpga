XlxV65EB    80a8    1880�0ΠĎ�����'�m�=&Τ/"6Av�����Έ#R��S�7P�t��t�A�s2ɝ�g��
簡ilOX�5Ix��J;�H��~,Y��Z�j9ߑa��Y����1�
>P��Fd+���C���d7��8��O�m��h%��w�-�5����$^y�7��&��dP��Wi��9��P�7���\Ǖ%�,���y�q�8�(��Fx)������x�t(�k 0{޽�t��V��	��S�&�����l�05~A��)����͌���oh����ZD��Ec�d�<��2��B��3�L2=t�BD;1�hU�^��F�5#s���)]���:���S�P���h�g��0��ʠ��p���ݯ��Y���8��hx�Ӭ�s'n䍤Buэlw��@Ҿ��.����on�2����o�ut�7��ͪ�$oO<�?���E�A1k|y �J=��������Y�������7J{��9g:�va=a��B��զz,���~��M�4p�L@*��SJG2�bA�⹄�a$?T}��^h\������g��:�!r��d�����c�GM�� �j�y��BY�F��{s��}���M`�!r��O 搅���G����K��g���XkI�y����	��G��!T=��bOې,�V�P������"��OD�^"%}��Й��N V�֐I�a3�_�n�	?w���VkS�"կu�T��7r�u-�%0��ϣd������n pMv�'����u9i�v�̮��,��M��e����������-v�EA���z�w��^�nge�}*?�D ���&����l7���G�f(��c�;���5~b �3�~�v5�%� :��gd��E��x[��gq6;ax��L^H��%�&>ΔJ��4�/�!�J
��P*��	����U}mL���2R�S͔���0R��&i�UȔx@p��Ѓ|�=��q��'Xx�B��I�]��X�c�q�����ET��]��+�rQ��IM�^D���fA�Ӷ��qφ�����}g����b�����G���<bvT���t����R�B~�+O1@F��x�~��lV�)z�,�U= �BE��i4~��cC���|����e����ضYwő7��3�q�8�bK��J$#�7�����6���J��,i9��)6D��Y"���i�����E[4JM���cc�+�j�pwM#��zB4��iu���5�:����Z�W�j�+N��)�H*y����^����)}��F��l���S�LWG�<���;�� ̚$LR@���W��*�)�2%�	�pG��-+��9j���^}�t~��N�,��U`OV�a[2Y#͐�1��F۫4�}��P�L͗d�k�(bvWGM$�o<��`Txk:?~x�h˯ �
�H@��<3����/�u�.��F���ojԍ,?���d?x$�Wu;@���D�>�8b�s� 9߈�9�e��i�_$��gN�����m^��yk�K�e�f��sY���_��z,�Hr"�7�$��dT�f#�UO_`�t�3��*pl�3R�]V>of��nG��<EB���Jaxf%ʖl7,]�;mmN�R��K�щ7z��w�F7������:��s��Eǩ�˛�u�����1�M#�L�<�\�6,���@�ժ3��Lo8�Rp1�|�x�%p =f�2r��ḁ����:�{�$c���y�Aۈ0�@V�$���-��=���-��$U��х��`46��}���`����8e��7@�Rݔ�J�֏dUO.pυo���L; vy��e�e#;Q��>���q�*%C��@�M�ӽ"e\[(��~��M�(wm�I�pF�\��&�HĎ��$B�,�z%m� ��T�<��N@8�"e��Z<N'��\|�Ƨ}�!�Lb(�}|��^N�`|��[��]E���A�Ϙ�	p*�jme䷦8��W|�]�%�#�&),_B�)���G��5�/�=*!�י�	���8Է�O2��-�z����M�&��a%b������U9�4����z}T~�wi��0��ً�?���d��D��7���c�s&?m4��S��6֘Q."q)��b�z�Z���x�}I&��ǲӊX�%��uv?���o�qG�z�t�ھ��ha)�ym��͈��P
N���\֞J�z��y�ï't^�R��7�ޓ"����Bҷ�iQ�� @������X0Bi�ݍ���y�/�q?��������u.�n����U�?�0�Y�Ou\P1��U*�R�W=b.��w9���4�h��`�O6�+u���e;�����-�ƃwӚH���}T��N�b�����Pa���=<�n:��E%J��ӗ����+�[V���0dة�~+:-�%�e$}݌�����3˅?t�׽'��$A�6�`����#j-��6�J��!L��<�z��'|�M�֘l.����V��,��4M@��K�&�bc�j���� ����)��Ж�ґPx]��!�(����q
 �;@��ɢ����h��� [�Dɾ����B�\�쥚��+O��xy�M'!�i����mY*�(�_l��x�nb�R��j����[��F%�Z����q5 �VG�fE�o����8��d0�<R�T��������}}��#��_���Zp�#lO�N�"�*��@�9��s�
i�Ի�q==]�" ˟Vc�јV���U��	f��7�vj�B<-���?�Ťـ��Г�=���Τ��d��)�L�4	�^�S�MR6�Oч��6؟2u�h�X�n�#�2W����H�Hv�1ǋxt�]�_�I���O���b⌾X�m�G���0�.��}�\�
QAـ�EE_��aK�ĵIn�����p�2|�
f�l�v���/_�����A��rd�k}Ck����{r���F&g5�oQ'���	�����[����z��S�ڋ=�u0����)~Cp��w���Ah�>�5=����<�b��,��6�5���Ƞ��P �C=CNv<�{{��:O{!�h毐�}Q����8��w��)�o�SOH��M nD֨C���݀yEUB��I���1z�mDC"�f���S4Ϫ�ĊWN-�زf�<gm��P��N&��'�Uu֬:b0%��U!�F

��J�$'A�"�npfɺFH�<��bDfm8�R���9��^o�y���]���C����3��po ���ter(���M]���oB��1�����A���0��	�*�\ʞ���a��0���@�0��G�-F�����t��s�if+��TdQ��%7��!�bI�\��ZG��b@�0FP �U�H��Ð_�J����]������J�i�]�'���	%�̬�gJ�q���Q���.�m� C��z�7{���1�wȘc-�'�'����N�x�bv������[r�o|}cz�u���f�ח	l�sG=�TR�����$�Q�Q$��'��w�+	���B�yjO.�ř]�׸�%�vM��9�8H6�x��{ϫO)�|B�ѓ�=�=p�)�I��ߥ���уMʥ��i���X�>x_D�X�^Jj��&��
_ٸ4��'g�qkL.Z �ơ�{i)&3�s��!ed_��ߙ���Z�s����ݗ�&�ϕ�^K���`������w4L�����@j+u�9��i")f�O�m^��D���Eb�&�Y4R)�Փ6��N=�)��������1�����c�At[�3 c�1��Z�S�Y��D���p��쒽>��%X>Ww�Z�OU�tI ����x0�٥w'�D�do�4�;̱8mc~�������</�ږ��Q4�Z#��&�u�t`vz�q���w&�e�g]���GU׎~k�I�h������L��%Ac��3���+\��#��}�Cŕ�m�:��섒�4�`�����k;z�~ &�M"�t�A�k�0�d�'.?ܒa�)77J��el�a�!7�d0�����J�+?N��^Cj14��S��]S���6�H�o~��� J�c1B���mY�cU�)��~�������3s��s�U�"v�8
�6���'DGD췳�wx��,x�+ِI��I걧�V�hK� vf⾞��Xu�L"5v� ����y_P
3�G��٫і���G�ȧ1�o�v�Li��9y�'�o��.��];^��j#�x�g]LJ:���\-9G1��.��sFmֽ��+aFmT��Hb���>�[1�saŠ�5���=Dw&��8�@f��P���y�o2�>�ЖK~Cv?�#>�iw�=��%N�y,�s4y����b��"Rdo�OMxs�U	0c�P�M�7��>��[�d�v ��~u��Y����8�t����|���>^@r°~)�[5��4��i=�t@��c���d�/8Mv?��ΰ���{���t���eͻu�K��F��4�?!h)�UӢQ�&��RҨW��v��lc��`�Ȭ��y�&ĭaw
<�&��2�)����/f����B�ؖ�
pv���?�fr-?��5���hu��R�X~�Z����&䝞~��F�r�/���@�>r?�&��ʵ�^(NP?�0և��h .ׄS�Π�iE�����u�3��KZ.���T��oJ�MR��j����`�Z(Ũ�Q��AЧ���<{��}� 2��z@|TP�,�Iί�	퐟V�?����/'7ݵ.��r��6��u�xw���
{OT�[��P���E��,X�>��`/óU?��!����<�Q8�������sb��?�`���NLƉ�����[�H��?Fl�|*�W���$���>W�Y7:�'Gt�vs֗k�B�N~mh��4]\u7+~��[�8H�Ml�(�#�X_ ,O��xWkU=:4�p3n;�Y�Y����_��;�k�� ������2�.!�bF�N��j�;]�ή��+h��&�y�ߞ���O���Q�b�%"�j�5rh�cm�©?5�삞'z�2d2�5��N�C�Ċ��o�ݴH��NE��6��/3F~�g���S��-��
y?2�ip�T�P�LG-��gqH��������+�x��!�
���]s��������n�
]6(sy҄�'����$��؇Ms;0ȍ  jf�U�ss$'EbJ���l��)Ȯʚ��%2���a#Z��x����8���ABm�J�t$F��u)�Ro�qb:Z�~֩L��� ���ˠ�l�t��y[��t��@!��-5��	`X�Dj;y���}���[��v�jw�F��l􌡖��A�"v�N�.i\,"(���j_6dD�ͷ]t�'�?������\ŵ*{ݍbRi��N�pQ�ٿʚS�^����0��<����|%�s-Y���F�����F2|De��DH�$.��v���jws���n�����������͈|+u��f�a��2�?�x[����zR�q)����T�G(����]C�����������g�౲i��uC�<�b�=FL�Ն^^w��9T���N5��hHۤQ�,�E�Ʃe7<BxBk+^��z��b��	�f��~q�V�"��Y���U�N�w�ƶ�T�ݪ�&��������:�F���W�7/+����Y�(���I���MR�/Y{�����r�.*�����y�-4�y���(�����t5=�罌]g�(�!RŚ9m�F��p|��]g'��q�8.rY��Ԗ�X��i �?,�eX��˭T&��N$�).���&�p��W�Y��̙p���p�҈
G�� ��B=&'{�Y�~&tW����5����e�䀌��_&rp��B�L'v=���3b���gk������=z䡯oM)�L �}�����m��G����_�?�i5Ff;/)Q�/�vvJ��hHX'�]z�+��1���������N�aV�\7��kh�N�k��r'�L��)B�4�4S55	xހ�^LD�28pf }���!"��#�RL	�E��Uj��>� FzΞ���t��WyS`9��;初�����8�gӇ]����{�Jo-���q�~m��Ii��	�����5�/��� �ղ��zp�^�ZꙪ�7l
e��E���%}/��C�Iq���n��K�
j	N��dR%�