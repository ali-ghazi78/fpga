XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����A�S�^���u�5'zs�yg�HRc����B�@���9M�����!�r��f��݂����X�z�>�iܘk�rV�oF,�yo�]}���%��	���t@;R<����<*�,�ܢ7rZ\�c��؊����J�a�7HW��wi�[3�|,?f�Zt
�PQ�#7b��dKj���F�M�BDi#�h"�ȢâӒv��	��ص=��eul�ʄ5Ű�j�R&7�7|x�G���bc�p���5S	�8X�\��o���L����]�n��_o����9ٖzXBU˕��e!����~�_Fh�/�Enz�UN�D�E�$?V��&�T3����.���'B��D��$T��r��5�w�f	Ά$��+��G��@�'6�BiӀ"paX�J���&<��C���>�	�� c�@��� '� tr�
"�a�v��SQV
��w��D�8��p���w���
�yQr���5 �6��d�2N��ƫbkT~��ߎͣ��d�w���˃$9@c��v<��s'��M媞��mHM�������G��[P���T@_�PHCѥ����JP�L�-Q!:Q��9�z]�bD��t�р[����2͔����w�&�乳ë�-�ʞR��=}�iW�ԙ�\�M��������M��2��O���[�����~�����̚~a� J%:�L��U�G���u�5�K�0�E�7=6���N5��9�+TD/���7\���+�s��nār��9N�H�=����M�p�qXlxVHYEB    fa00    3300��ZCUj�iUIkHjt����쯣�(>H6�[+s��Qʰj_���G�2W��״7�E���dJeG��k�5#[ʿªݞ'Y	w/]�e��������ԇC�C���ŭ\�1���tt�J7����Iu��*�J�p��)
�\����d���a���f:S� ��=�}Vb��~��#!�Gg}�#\6�|�[vV�A.���x�L�r��3`����`����HG��>)��T��kn��}��&��T�,܀*�SG�նa�\>�����2�N����ĠpC�FS��Z���o����q[ʹ"���QV�U���>G�+���-��P�wOd��'��Kz��1S�o��u��M��£\��Id�� *hE���0�Hq`����������Q����X�y�>����.HNq��O��D�RzȮ�h�"Y�W�y���?�T���ǣ�ALt�v��7�|�a~�K�C!~c�JyvE:���ut�P�O���uzr�,��(�䙜)64i�_��+���e�7hy�P��BQ���=y�^�	-ى��W�9��^b�%:5A��g�9OSΐ輒|M
j.�v~yC{1�D�^{f�]U���A	�ft;�ѭ�>��*�j\�%�D�ab}ΰ��-�1��{Rz���ҁ�7��9%��m�]��{-����d\�/y���+�M}�s���	�z[. ��0�!�ޟ͝w(wF~�,﻿R���mDR�@x~'L}����m���M��e��p�����8��@��_�X[�붠� 1����nZ�%��g��s��,���i��ޮyW����oC��'h�Zk��how���.�*�NX��iг��>��s���F����kY�y�gj�˛hj�ϸ�ꩴ��+���ɕ�S�ț���n1��}'[7!�Ϝk�lqd��ܓ�}��M�w��=�%6��|���ϡ[cṽ���� ����H%���Ng)aŘ���
�A�c����'4��O�V�����V�����}@╻ӆ�0ˮPaFkk��\k����գ`������t�����BB"��6M1�@.8�D�k��\�궕����v6��e���yE*.�v*�ƫ��|)�W��p����j�9�D*�MC?�9m��<�S�	p�P<���ޘ[qM��� A���ck=��r,_���(J�U�ZP��
��;��/.\%�(\N�YAxEs���ͥI�ۗJH:���!<�.9+,��`��)J��z!�+�lC��;��x����]���F$4��ܟ�Gݍ	`I��bX
�"���<?�;ћ�����]q�殑��N��|Z�v���J���iBU��MQ�q��(&���?��e=����!��"J�U�&�.��~�8�P�5��%��@����]���E��|Dm_-�y�]����S��_|K^M/�v��f3(��(�Gp��J9�_�Q,$���tA�P�����;h���~�q�]�s��l��i>�U�}'lZ�at����Ê.������k!L�,�UJӯC8��Zݿ�A?���w��T����� ��Gr��Ms�Q]����2e�-d4:~Zݛ<삻�S��J����9���S~�X|�Dt_{���r�9��\)=�`�T�l�r�V��(�0�5ğ��]�R�"����l60����n��7�ߘ�"JW��a�t���0���sx��5���?�R�L��|�����R1t^p��cݚG�o�> B��g1<W_�I帼���D����8L?�O^	��,E��8(���=�8�����ǩ�qR���K�яH)��lN �ǭE�^���6��:�M�I����+}r�:KG\qsS�M����3Q>{|�7�� �
�i�*�/l=�)�k��u�a�冫�,A��Q(�s���<S��Zz�q}�a�h��e�R��Q�$>F*���N�@*A-�N�d�ə&c��.�f��/< ��0��������A�'��̞w�a��c�x#Ov�5�R�kO�oiB��|�B m"/
�zu%!��x痽qU�si�d�Y<k��%.�'S7��� �K��"�|�w@~��ku؝4�v���.C��6��	+K¬�ف�\Ô.*�g�gB��=��p�_x,�(�m>R��������5?��(XV��ӫlο����2���\g%�Ц< ���h��q.����Լ�^�@��2M�=��/�lƾ��-:��V�=ށ1�Y�򴼄���̸��6N�A�v͖m��<:��혆�O��ҽs�}\�n�[l~ ��	9�7���~~�t�8>��~�	��yU�t���S������!�@�2,k!p�ޅ�a������σcb�=�EV���u������L{p�@�f�>����k�����!K8������(�l�n�:�N�����J')�cɞ��	R�u7��K4��'�nI������IW��/(B����K#���ziU�OdB��<m�^�6[�qK�UH�A��@(d����`�N�Mʫfs<c��8�R�P��r��i����W�Q������_|3�:#fQ����_(���,��p2��#�"��]��̆Hf��NC�)���|Q/�y�H�+蔢�L%��ݢ�yj:(�&�f��m�6��r+�#��o5�|i@A�Xo�i��.ߥb��%�9oZ!jQ⸺X���cQr��U�Ʒf��	�^6RIܻ�"��������rbR�D4�G����r����u��?�x�]G����h��j���jHQ�.���B�%)zs�h�;-_��0+q}񎜍*~i����A@N���4a���j�]>��b�(��dX�,,��J�,�B��:���o�iq��?��Eoޤ�-�����ju�nਡ��9DS���M{m�|��^b��G��Y��
[�П\1z�$�K4U�'�[����z�f�ԃU�� }��cit�ǫ\.NZ�XL���¬��5�&�|��h�M	���X��\ފ�FB3߾fN�nn����H�eM7���u�� :#�g��:R9ts���U����<�C�u ��z��Ȗ6� F�(���j7dNs{��5A�fJ�
T����+]J����{'c��,�#{�����'�w���J7���g�-���{����eAK�F�e<�*�$"a��H"�_��۴������f�H��n�d8q��B�*�O���������~�S�!MI�SGH�"���V��
1b�^$��=�c�5`}~
v�L���c�QNɳ����	3)iΉ�h��:<=�@��w�3_�=�AXMJ��7 ���	��Ux%��i���,�6�����O9�quB���DL."� zN��=�v[pRU�9j�l�����b�قM4v�)���ރ����:@�Ȧ�I���My��cl��c������L;фO%a[�8��g!�!���ᵞ&d�Xy�̑ Bq���nh�Mb_�nq����y3"J\��bLE�
�����-Ԉ4r�5���wG�C(�b�+w.x�����c�����$>v�*VV|q�ǩ���݃l�P���(a��&�}^L��4}����DK�\��y��Rכ{� pl9:�f���K�?�M�8`p�m$���v�Ġ�c�" ���P�%�}�h>��{#���!��ܲǴ�P@��w�y����� ��򭕝/"�����͂o
�.د�|�*.;����C�ۈ����}X�HA���3��`��ɽ�FV���ʓ�u~]���j\v�I�7�>�/����-�lz�
�Oc!��d���8K�D|a�������m�v�l���y�����J��Ҋ�\[�:��'��,��_l���Av�/z�)���(�bOm���	����|���lL�!��	�g[\21�H�/�Q��'#�R��&�̽��ҩ��Ig��h6�N�� ���s$��?���?v
I?GD�B*���{f��u�	��w�A�WO'�q���;��n��U٬��=2O�t��t*�)���:�J�_wF��}�b89�Z:삑���ó$,㟘ԥ��F�ݮ7�֧Qf�r[6KaA��$��g�Q�Zzp�����1�cS6�0�Ҡp�i�B�rãH�����D]����BY	�	V1(�t_�>��M��HA� ���ɡ��A����lT:U�a9s��Ek".L����6����a8]��4[�������u�v"��8�osD�[)��.4E�~� r��l}(��o��-�6#/)�$v���)y�eoѪ���BW�j�����?*Y�2dU�|S��-׸�Ğo���H�u����'�^�Ė���hz1:�J����xAl��+�ɟВ�<ٰ8�q ��`����B�YqN2�-hxFm�8��f~�J֌f܏�Ғ,ZN`��B���Ք�4�hK?��6<�2WI����h��?�	\#�$D�'��"?/gL�jm��MDG.R�F��
��3�9t?�Z���r��eA�pZ�,�E�Sl��(tY���4���PJ��Ob�P�5��"1�ӭ�͖��34EQk���@�������=��5�wJ&���Nt�u����x$�񊌡R'�D��ܻQ����k�WN��H�B���$Z��X�C��e�8�Y�l���t^t��D�6s��5'V푱!v��;�.8(���&W$29ˈ�o��H��P;]��H��W�(���W��H̖�=pu]��د�|�R�cEp�#��Uk`��<-IϪ7b�r1���\���N�e[��2�e\����FԪ�ҧ}��GO$Q��/.�J��N܄!�K�'�SJ�^>�S�l)�^`�ʱD����`E�
t���E������q���_:P5�Q<Kک&�!]5\i��i*���J��������	L�2�XLk��)�<���<�9��,Gy*��T����q�2h�f�������^D���zsĝ%م�$�z���>��x���	�2��R6=d�ժ���@�cqMoHNa�L7d}�[�-�9��Z�f,Gk� {�ߵӃ��8�@��Z�W���.��U�G�N�p���])wϯ�d��[̯���>{�A��N�{K(��C�ʳ������:1�r�8!�A(פ��.����7�r�� �=�`]���җ�Zq.�6��,���TF��$�` ���8�	bt7����WW������:��*�UL��@���|7�\�tZc�Jm�5�-O`�^-�� ��쵃~~�i��c>�W���7�pv��l�k%�>��5�ԳH�dtx4��Y�|ed�X� g��9��/V�GH��1yg0ճ`��yV�L���x��������ņ�,:D�'�QZk�NfZN(o��~�ÈFexO����z4�
��1��NQw��&��.�X��Kt\�0�0�X�*�J�G펟E���=��<�pB_�\O�3��.�F!��kP{CZNf"��|:�P.�ǔ��p��;0ÚϨZl@f�!�_��F��z�@'��<Zb������V��X�'������;9ɪR�|!�Q� )�����(L�bQ��iW�0 �j���E���$HC��n�t�p;Q�,�Q��5��P�g�q'$�~���*��ڝģHm��7���l������ϊ��坰r�Ai�J��#��k��6���:A����譩�z�L�d���^ً�S]^�8V����1�^�ζX�hx��h5��ٲ-*������L7�?I��x5fmz��Dn9�j�����pvW���/��w���;������lr����r���%;�>��_��ـ-�'d}L&P��_Uw�<��Tώ�NT�Q�D쾸s,�9(X���y�@�e��~\g7c�_pD%���Eƒ��j���Hݲ��FR~���v�x_��$��x> c{�8,�o�?�T9�K
 ת*Mn�������ÿ0�V��O�8o+hmA����	ٖ�M��t~#Qd��ł>�&!��1�h��h8>��@�=fС�>Β�����d w�Wө`�h6X#��V	{!��P��7$-�T����σ)Wl@XP��iP�-5���5�PJQ�/F�aNH�����V1������/5|&��My��&��êsS�q��K+d^��T}�������V�=��n�:������%�� 4��r����ԃ�j���;ڝ����ʩ��	��*�Ҍ�1���d�e�9�k�MO_���e�tOp�(D�Rri"�{�b���b���<�d�m1�7���[O�_���G�^c !3������m^Op��̟�Ҙ��d�t2f��|��o��E�x��m�<�#�j~N����Տ�	�1 ���Z�,`52K�';�,��<���0���4gr=����q�>���Q��)�:��ae�N���&5�{�����cKKZ1�6�q<�/��\E@��n�`��@V�r��ɰt�Kr�h�b>�+@�%��yR���N���ۮ�`!����F"� �h���o�dG�IΤ~�����Tlʛ��a5G��f�,�8��$��S
r���)�C���C�����︉�A��
B����[d��]`-�쫨�q�'�.�
_g}�繊aP��~���K�=Ƙr�V�䪇a��`���c*��O�O������hKV)��d�OX�**#��2�\�P[�~�mH�]ɨ���G��P���I�hQ��=��(�|	���>vXP0��
��&ʼ4��b|�M=��6�A������8�M�_7���!���q���b @\�=>�vhA��ܨ���}�
ـ�99�r�,��DѸ�u��Nc�\X���e�C"h�� tB�#{N>,3�/�����V!���ȱ��9�� h��x�X� I�$�qsFnDE�Ri�<\��� %���~���U>�3��&�i5l%mxǪ���$�����l��H1�jF`�6��1a�����G�*:,j��������iNfWo�8��]���� ��+����0�^Lss�i�}>�J�/)��F��)E�ތW��[����Q*&z����4u"�v�Q	�7�g��k	N�:�*���q����g�s�c6߀X�*�o1�Q�����f�ZV ¢z`�WVt^���_�$��.���&و�UhEax�xUS��7
DT�]�c��=�v��A\0����ܼz�I���\��P���r���v|{�B�k
��$�_��P2�ű
C�LXē���@3���"��3Yg�!��DW�pl��0��Wi��Pn�g�˭�s$N������ˎv�T\��v�TC�����?,�Ԁeڏ����2���L��Q�yE��Z�l�i�6]�$�0$Eg���M���
�P}f�?O�a�|�w<;���v:�T-r2�"Z�=s&֊>������"�kP��s7]'�݂�S�~��U���D���� D�±#����E��JP��Cr���3�n���)����t}&S)�(�s.�1qO���#! |i9����*����T`ǃ�áS�NƂS���%�4�bU�Y�{ɾ���?KSn���T��A~�L]J'������{���8mL�?|D$����t�h��h�Z��!S}�+��|�D*��/���Nl=S�WX5��VQ�(��"��s}x��u������홧g���tLG[��}~Բ/ۦ�'19�B���׼��������^���y`dQ�o�P�es+�W�O��J�Ћ�%-��.�ز¥b��{��	 ��>��>~2;�)d^'�,в���>3`�yo �6LG`@��v%h�*��+�5���ޯ.F'�ۣ�޽�>fT�=D����QLxZ)�/���E�`��DƟF�:��yu<��������u|2��q�#�t�$�%�mF�2LotHd݇ow�\�mG�_;��V���Y���q���һ�(=0F��B�yR�HI\S�H��=�����A޴�N5��Ҭ=��`�#�^�W���,Nrhy�������7�LF��b1�r�%�b9T������"�R������d��k�HѸYa���|�}xF�ʷ(n%e��V���b�H����й�Z���mF�o���۷$u! =�L��Z5���Τ�*˳�v����3tՎ��­	h<K��L&ھ~yUE����~���:6�Bk_zN�=���w}�'z��ͦJ�X�r�t^p���#5��~pTPb�. |�NRY�q�C �lf��JԲB콉f��Z�S;rB�˗GCe���}Y~�{���i��e��8��̻�n�K�/b0-�'�ϐy������f��8������ى��&3;��|9�W�{՟�\�Y,Y�"|��`��6ʀ�޴�!ܹǫ��V��3�iM���wcQ�c՜�ӘU��߻~��4[]tT�3�&o��D�X9��S�\XV�I��P@�~5a~�gx|��!�z�����5����=S�}j�g�g��X���ٺ ��	"e�#~�O�I��a�!y���zT	�ߏ���U����s5����jYo+Ź6o~$�9NW�d������t<��JJ�_��@l@H����a����� ���w�AM�g(|&�V�w��V�^sYe����#<�b,U��n��,~�d =��?��;̦��ȓ��Y<�kҋ觽�=�h��۩�J�X;y�Nj�G�����9��#>H�|I�{X����s�?���~�Jփ���F��AC<m�K��5�K�uf5�5g���g��.dM_���P��G�ox�hT�a4B8)Om�?��V��|�@�%�e\��vu�5h#���F��)L��䗍w�p�P�#���9���B�P�&���6�E��lzVH�.Qc�$W ��~Q�U3��0��yasWa0_+U>b�SoF�Ql����,8����W8�J�&�
^�w
 �����	a3"��E�N��S�5����>���� ��Z;�o��gm��m�����ׯa8��Qn�)V�B��l��&�-P�n�Mx7�];��I�������0����H(��-�%x�~r�n�Ŀ��� �\�v�����:�@�C�m��gZ`���Y�4���pOIfQ�LѢ叙_�������B�G(�fr�o��`h���5=p� {�ݾg��ワ�d��أ�2w�8
k;�og���UV��F�s���H�ߋw�qY�;]-,�mG枡œ�[b?y�B����
Mv?�W.fK�6W��%����vl����Bș���DH�^���G;Y��Y������S�'��� � ��~٦q5��������ۂi'�&�a���]o�����(v�Zt�zZ;�#ʻ &IN,��s6�C�9��b����/_nܱ�pb�y���<��U�л9��1O�x"O����(b�@����>7	���q�a�����m�aU�A�z۞o-˅�߇�nԚ�G�N��m� 	j��J�Q��7��S�	�����kZ�STM����$<��xT�.�"#`~Q*2�tMÐ��x0�dq��B���J}P�F#J�&l�Қv�!{8i�O��k�1G��J ���XNO�p�Nm|������=3�0�bog�ɓ�����AJ����j���,!)G��[��2����Y=�z��"�,ׄ�e���e���<s�R� ���x�-����&��f�ţw���})@�T�-"�U �u>V�m���uK:�R�'K������?K�/>���+�&�9q�R���Ͳ�7]�m���,П,�˞>N'KB�S����B���Tt��AΚR��b̔�T��+�H�o�A�63�� �p��S�}f�e�R��y�2+�s@"Y��}��	�݊��8��C4
?�Kt��##�S�i�ڼ��36�;�_ןi˼��p`�j� ��4��f	e@�vŦ֞|^��� �y�+��珽a�W�}���[��~�I$�wB����N[Bm%�1�V��
i�h3�?&�k�2�M*J!��p4�_�*W���|���;��'C�G\կ�<1i�D�7B��'�KS�m��t2�����l��A�4��ׂ�w�<y{��{��5�N�+�69�KI�Zt���87��V����]�	0&��~[�RV����WD����(�ƶ�ȱ��̓p��+5���>)��C����������C=�sa�����rO)���Ͷ��G�`\��ab�G�&��^b�Վ�x��9���� ��f�\��<U���B,pE	����>����2���r�'d�{��<:��޲��Csk�\P�\�k8��Uw$�"�J�R���sY�ވ3R7���x1	���wն('�(�9|�*}�ظ�S�@���g�X�M«�xha��S@����1����~M�����Y[w��9��qH��pv	���Upeޥ`y	4t���u2�����r��~�L56�%z5��R��(i�Ω����C��;���c��bfZ+��ʊ�q�M��`�C�cHYh��r��h�4�!�6���Zu���nN��D8�����ϳ���YI���1���{��U�v�[f�)���r|Ȁ�MR<����ͮ�(�PVo�"�b�+�U!(����5K��9n`C�M)\OxZؓ�M�$�@/��9����(�+1�!
��@���=����/�s�
7ñ0��6��S��0g
�:�-�!0����)eM��B��U����y>�J�>��cy���J����$$m���Ǫ�P��B�۝���̖E��6M�ܞ9�H��|�B���9�c����}���x���ת�uYP�}>�mVG�S�ԳO�t�[�����[���g��d�	w"w�p��:��vq�n�6u��a��V�|���V#n*��j��΄��7�a�@��'>NP���N��/
�j�i�s��-�iW�q4R4��{��)�>�-tf�3���i��&�$̭&�;H�ع&��#�$=��i�ug��/X�z���)�,�ya�蕧.���*.��n�q��#]a]���@@F�l��:'\��f� 5��}5�&�Ƚ�9]�01޸9�(��lX��/���#+\�7��U�w��],���%�o���BR=ɨ�	��}��P���f&����	]��V�٥�8�m��C����>�;ʜ��a�k�䦙?�b^sײro�΋�6�ؿ�]>��5���ʷ��	�[�|sBKno8k���W<i�~���52K�T�[�5�L�v�n��÷�-_<���,
!2�I��:�u���[�j�d�7ͬ(��U�����}��\~��#5�5�W%� ��r�S�F��wm�g�}w��\�6���$����"�Fw�7`!�x=�����JKs�l*�m���I>�*=��$ɸ�Ag�{��bڱ�R=�:��P�?�j��G\��s2��<�s��Z�ץ����n���#<���}�r��Fx��݅���EwlE$�����Z�*�n�c��N�:L��%�+����*G=s���h��?T���r�+I^of̙gxZ.I/e꫅��d�3��m����B!1Ќ�tA�2�$�c�S���p(�/L4ND��C�h�����Wq��3�ٶ�y�����A��,�B ��ݛgI}����-���Ӵ���ZT���)ں����w�Q�jbBOF�(�9�NV��E���C��.�=;2K���O�A��Fx#6߼I�.J����k��8tq�Ψ\���p.湉GLS��2�~ݛ�������%;�;���FQ�`�>޴�"݂F��E�t%)ϔ%�p�rKqfS�|�����]�#`Ǩz���Ђ+�+��r_�v��o��l�G���b��;S9~���f �?r��GB�����n����;�w9mnsRJZ�I�k�2�kL"=	
3P-a��~�Ͻ���dr��xw!�ͻⶀ~�]��73v�����U�v�u���
gQ�%JdނW��U~�6:�>k|�/��Se�^��p2�>0�6>��!��IS/1fY{nn�=�pj�QxK�ǚo UL;��#! GD��~'g�l���9��JK�]��s�q�,u'�}��I�����Φ�jVr�dj3YE)47�EC�Ρ�d[0`���\�'��\��Ի�C�)tTܴ�[$1�Z��Q���2�7Smq}��w�kRi�	���}&M(�dM1�4pۣǒ�6B	0g�E�����ac8���h�C?����ġ��O<S��^:b>�1 k��BB���$���5�[y@7w�A^�,C[B�3�~��,���~�l>�V�+���GH(��w�p�Q�K���h\�cN�+��}֮o�)�����MH��P��4Y���W�؏�=zD�t�,�=�7u�����"tۋM���N�Ci�"��0,w�0-		�%���t1.x�Wz���&Ei����ꀱA�Z�1�z{�Jhf�v��3y���~��C�T��7C򸡎.��.�*o�#����xtZ-)#���G�ϵ2.͚`sJ��0��=؝�y������Xd�����J�x8�*�#?��[�dX	 �0��M���թ~=�D���,vS56Yl$`����-A��c������dUQ4��^+b����2l�O�WmdQKo'qy��Yh�I���>�W��U^P���z��ݡ�cݟ�"Y�����5_g�'c��3�y�a�̴�a���݄^fP���UX{ꧣ�.�s�*����5�6�6�*���\|�O?��Z�;�`:QG�`DPy�p���o��za���W{(�=�?_ο�Z8�S����`��3g&�R1�	pEr`
V|�t�j3%�q���XlxVHYEB    6855    14f0Aᝦ8K������s���6�Oi �� �aP�������`�����H��΃�:��I�ݢ{K��u>���Ia@*{u[pm�Ŧ���	4��㬤DQS��X>H~A�������}]�����t�Kja���9��Г�h�!�ۡ�(0���x�y��H0�� �����(E���H�������E,N`~�ɟo bJ;d��������<O<Z��So�8p�<u�f������i��,q�p"����C�A�ݛbì�av��_˖�IL6L�ݪ���n��8Y�P4��ŖҊ�U��u�jV��v# i5ѻ,!.��!����9];?��u�!�3T2�'�,/��R��삥2�\3V>�$kV���.�]��,Ls���GF �W ��z���{8CKw�D�^Gɋ����Y%�3凕�!o����A��@�h\������:�>`�ٵ!�(��lZ���E�~3=�`M�q�DH�EP>8� P;�����ھ<̩���(����S�]ϛ����
798���5̞�6����2 �!��G3%4*-���q���`�Ԧs�C������@Dn�?�*��X��=��A:��d4/�K��x+��!ӳf�%^>k���?$?M�����Hhh	%�񒸖s��%&�}��s�σ�vP�D�:��s`����+6��}L؟����б͹�r���}��x1�X�4*��.�vqm��D��7T��2������/YdJ	8T�ˏ�^���W��6ՓL�w>��[%�4��t?|�@qrx��<l��*a����b���}�1�.r:�P���OV�<1���^5�u��P��	"�T�U�z ��a�8�I����Lb�W���+Ǟ���e��{v�"�V��,ƓO8}�tߥ��'�(���5��w�a��a��XI�����������^��D��=Ҽ�k�hR�q8�Ōdz��v�W�HD�y��I��VQ���y5];���Um�R0��՜t+ǣe����*�i�谌m�P��, ��n������aǀTlH�]8>n@F���-�f �-'�utv~�r�8T4P��K�{��X������+=3��~1{�+����}m��j\D�kޝ�m��{D�{��r����B`ʍ���� �|(Z9_�]�Bc�[�G�I�ZTO�����4�W��1��/�M���A���#Ά��k����'�!�$[�uZ��Oh�1['=^�\��6���*��W���L��	IN-p�{���7{ �RJ#|*d3����SZ�M�*���4�K�4�ɘ�-۸�PuT7�1|��'tׇ,T`?��'�6���ܖ�'�<~eN8V�
x ���,=�-�{1���J����|�@��-�I���*�
t�ZL�;�E�ؒs�aa?��EN&�D2Dx����ώ:ָb����=���,x���T�P֐��҂?�g��n,��q��ʒ�)���Vb�*3�2���)g�w�<^�I�d�M�1�:'x��!#η�NEy�z���D�a*	1��uF����[���e/E��R XwO�=s�[�a�,W#!b�q�6��=��b���#ͥ�,�Z;p�Ϸ�^c�d�A�Y+˝�ܯ�i�+���kjtm��m��9!n%��s�t�V;T��(k���Ԇ�R!�5������H��9
���'�F��A��{q�ܛ���=�o|M�KA.���"�G�]w9���[��/�9��'��<�+L�c����/�5+;��V<���t���:f�3P� �.�/�����x���0<.h����Y�iQQ���s�t9�4��4D�� "��l<a,�n׫j��S&���9h�_JfhU!���f�d?�������"��ՄE�;,zR�tx�/Y8mM1T�`Zo���^D��`��E#{��PJ�wҝ�+p�S�z���K�=�҆��i���h�nRҎ�B��E�ب����٢�4*^W���Y��8����8wQ���f(ù n�W��B���Š�x����L���
Ye�U���E;3^2<�J-��,Y�π?&o۾��� �?��B��FV%A����� ��h�}@&�0�����w��<V��u[%�ܓ���|�*VP�E%��P�mU�<��S#m���i���@�;�즅� ������<g�s�}�K���r�b(9^��������{l ޒ���VIov)l����\S2SW��J �7x�Yi���΍���?����Y��|���P+���gj��=b�h�$C+@�`ԓ*�H� ��N�ȩO�
�bKz1ȕA'i��Β��W�\�q��s�AG��Xޖ[��a��9�D��3g�_o�b%[��i
,f7K�b�0U��k�a�$��
H�8��L�x86�M#{���K�ILz�8�˞�n�
j�A�}�_]��d�/N���ּ�x�:�^�p���D�r}�(�^���Y��W��'7��� *=�Τm�a�|�-��*:�Sz5�:ke�ēx�(79yj*R�\�[;�\p����K��:2�>e�ACY]���A$dC���%�����gfj`wZo'χ��іA�XA΢0]t�4�6��E����\�9�j��@�e=%6�U��H�Rr�J���u�Y��b�B���2����.��L��Vr#Y��{�U$';R�;<ڊn�TDL��pH�=1$O��m�*#��]+4��͐�yB�j:�X6��,u�&��ݹ�����2�]AE%&�U��9:�z5(����������^���6Ԥ��t�N)7Jo&�����#*~�fdi���k���#�<�P9���As�p�,��S(P��KE�X��6b��4FW��V��kU	���g�J�T���΂!e;W6�EӡK�t˦
���'���l
D��8.Q�:�X$6���v�A��\�6 "Z~w]����Z��<�\l.�yQ�d����ȓ��@���g�_Z��,��������br����8\�a�N3P�aO?��i�A�U$j3�Q�'l6��2ɀ|F#����oiW0i@��eQ��1/L����e����i:O�#�9��l	��RA��H��t�}�̔iS�W�c`���K�BI�����Q$(��m��-�X,����Tn���w��kS�W}�חȆ�������q_�-]��ù����Ԋ��wb�n��:�7<��R� n�L�s�D/h&�s:�r��ё�N.a�Ɍ#k�G`c�ܮ1�<�[W)13w�<�Aî��S*�̭P�+ً�A�	�E� �Ϧ�79~�=^e0q���"h���x�R�ď@�]�i�0ᑟ?����#n͠�m�1��З[B3;��CĂ��%������ȵ	�X������pΜcS��:�\���|Z�:�:X�!�M�vn�(�\�s��Ȭ���I�""�\�c�Ѯ���S�>od �Q���@Ud��H������Ǆ�2m���ȟ��e�1<9���	Tk��P�_$5M���_݌N��LM����(��Aq��yQ���ɡ���L����V�(Fk<���������M�/�'�:�J��;P�C��v��.���[(�+�Q5.�[E����AFm�!�����L�ލy� ��k�t�is���{����y��?.�����.�8���W�QR�\�b��m��l���N�����
e'gP}r����� �\VN���Q�q�9�x!��9�H�s�Y��.���>Yw{逖�[��]"bf,q������A)�e"��`��au����l'�����żֲ��X$Q��,1��7�;��v:X	p��1�_�y_���؆�E�s�������7�9�`F�n��L�$p��JÞ�1ic��F�b�($Wj�R���uٽ�\���,��{����pwY�$c�l������ݷ��fw�<�g&�s��dBDd��<�=��;�ǵ�9�t)*֖�4s��� q�qL7��&�\ Cf�?8i݇/������zj�@
@��ؚJ�F`hD1�ѧn}�Pc�P�+UHn/?����u��G``c��W�����eN[d��C���%���@�"ß�:�<�0��'��I\�������K��|.Q�֞���"�Y�~�\z��8��^�l�ɢ�޲p�y$]�:�rz�f���k�������Y��C���!�(g��J��V�Yt$��E�!�w�8n+���{a���t�A䎗�{�XUɡ�7~}��i+��n�n
�j�7,�p�H�6�L J����յn��Y,?E�N� X�^��8Cg��Ϟ��C���1�A��i�uד��]�dM�`����/�Y3���pc�I��ÍX�� +BQ6�D%0���byl�'����n�^Q���o�����P~^!��?�����'�H�p�����.W"�*A<��%@���TeD�oB�ǒ�=O�2��rxI豕a�8:|(d���6.F�&��:���prv?��k�'oP���Ԓ��������g&�������o,���ƀ-ɧ#R̄x16��/���z���m��?t�����>�d�n��"�b���8�J�v"T���u�CX�!�v/�LU�+2s*��}o�/0�S�߃��w7૓���e�bN���1
��^��?�P��RƉW����R���9�zW��%΃���d��%)oM[=6�V�q�m���+~�(տ����&��ta�&m���x�1=q�V�ЧBc+%�����O��:��N~���A�B��~�g�H�x��X8x�$S|e����ݚEHD;O~$J��t4j��t�e��'t�Ϩ�GM*M�q������<De��pe�>�MQ���.��MD:�_��+H��	���`du�F�猑uz0~<�ԑ>�Q��2��8�T=�+�-�1���DZcu���)Jz��9�,d��L҉��M�������A`hT�P��H��ե�2����N�V��KY��hl��jJL�C��쀍���"�|"���Ei�<�r�1�:0��3'��fm�{�{�C[s�`k�|�c�[b<�s�'2��Nr%����@{�`5��{�c�Ԓ��/��*���(ewPX���%C��2���~b�.6�=L+sle@���|tK�C�s�3�w0�b��y[mv��(��	�5�4Os����"$/�YԞWюU$��;��[�{�*o\O�AЙ�h�N�#���A��Spc�Ͻ�ga\�ۻ�<L�����;t՗�62�b/W�L��_���m�XenU��,G