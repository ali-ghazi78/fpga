XlxV65EB    5289    11c0��?�Ƽ�*q��R��� 3`P'z>7Q&���nT�8�,�(�4ksC�T�ԣ 3V@n`0 �b���CS۾Z</�(6="c�X&��a����믔a���I���qkќ {L�7���,l;i���ITݒP����dw'4g|ڠ�ne�����]K�|ϛ[	G�Ȍ�S��-�fԅ#(���V����%|���1g^f,x���ώ�Qs���n��Ij0����Y��c�I�58�8��&�}���6G�V���yF&X)�Y��4\�0��T�
��ݟܚ��#�����=���DqPR����8i������p�ܷN������֪�P��b�bS3��q�������`���<>N~P8m`��*��惋�8D���r�� t�O����)�P)�7K�D��S��!��K�5P\<ЙWT�7UE���y5�I6����2�0*L��-d�m��t�; ~�{il9����W]�(ӛ!� �\3��3��.��1�����
�wm���0�ƣ�E��
ڿ� ;��7JE�׉X1�\���bm������g("�5(�d{)4Y��n��+�;���rl�/S�^��OJ��6�9�>�t��J^ź\b��=;��]�������?�尃�7��� '}�T�ݧ�`ͩ�k+�t%.��T�< ���}�p"mt������ߵi�߾��S'�A�<�]�ֽ�5(��-n߯��8i\" ��a)ˣc�H�r�KU�8[�w2+��A'��Vׄ@"��7Y9-��%����2z��z�S�̚��>>���m2�RVd��"5�Gp�L.]n(�<1���'3;y���pa�\�;�Б��s�Y�1|5������;�c�}Y�4P9�����y�5������u� �nt��;Z!�އ!��zMN��1�e����U���w�]��U��� �yYW%�����ERu�4�� Y9uP��n|84gQ��>/��k���Ę@�!�1&'6�X��㹂�gH��D����5����{��ot�Jlpv�ҥӫ����X�"A"Y�.�}�,ev���2�t�̏{Z��u���.�BB���v=;�S��V$o-�������X�@t�	���7̋*;��Æ3WrKFb�׆r���[_z���J����fzm�C�F�����H�.�Y�{�հ{ER�y�C{#&��>��9����!S��d�q���Ù��s%�+N7��3)M\���$�����g���M�`�>�:R��\���𻥒��V|	�+���y|F�OF9�	̣���c|��kK���:���U�F:q��;�����6�k�1O+9f��߳�+
p�z��v��c��I+	�t�IpY|�V1�1#�)A�3��xh�N�%OoG���p��&�^��x0 �/���G��|^T��	�J�#�4a��X��^�@����1)k�-�]�nҶ��B� 9
>���匷kJ���	� ���D���I��s��u��Q���R+2�No�Rm���.���W\��3Ű�X1Sf��X�M��Xa9�ݰ�Z����Q�W����M?�}���&&�Y���zk�Oc?>1Dv��M_Zd;i�<����=뿅K��Y�J#Q�� �NdШ��T�� ����r�}�Q`����M#��ʕ'N甪i�&�u�;��Hc9�8̨>3�״v`����S;u�!��-帎k�*R\�?�E��!;]b�)�=+�������"���cH2rB�SY�SQ��+rZ��4�t�MAAm�΢�{�3���S;�jpe����b�h��2�?�%b�q3qX^��X��jtd|)"0'�7�<F*�yA�/���Ġ#�e��$r�;-{2������^�C1k���w�p�P�tq��mX7~������j"Ƥ ���L�������N&�n��XB�����F j��� /��u�t7�����%���(����B�O��8��[v�W���.�a�%���8��]�i��P<\I��пX(na��!pL�>l*���*@�W�z����WQL���_��p��]?�\���G+���*�)�o�]Rh�c@���ro��>�#seܺ��s�	=��yL�FK��ӛU�
�X𮰎E�)Fd�)�,9�5��i�_�2o���#M\%D#�j��Ê�@�x6]D�{P�X��C�`����L-�P���*��P[�_���� ���r.��m�9z�x�	�^򖨆�`1��q��q���v�!DDPC�30��HG�?C�)7�ﻳ~B�M�O[�֚E�K�!�N��	���~��7�US	�G�:֋���xa��$��|��F�R�
�Yl�S��6s�V}��Ր�@'=O��Ĥ&�lw������D�y����=#��|=9/̰}%�9fX�E<nzvv�w�8t�~dg�8Q�}%;��]���	fvh�R-ǈ��g�&�윘pv�����Q:��*�?bC+��*l����\��rIʦ��g�`^Ί��NqG�u}1>�k-��FN���w�JMK;i�ĝ?h����Z���k����uj�QE�#�C�U�˼�2
_�g�a�p[䰒.��e���5��$�$O�QN�Ӝ^����1�	�����/T�o���������B�����B���졹7UB��8�U����l�Վ�bx>���L��s{�.�:�53܁���>�1��7�e��}�:1v$)������4�0�s|�!�����={����fK���3�j�?���u�J��N�Y�>7���Pf�qÿPִ(���}WN���ա�g K�Y-����������K�_y�ͳ���i�{	����G��q�����ɸ&~��Ec�.��mFؔP��A�4��iLx�x��eۇ�.-C�ŗI��\?M5Z���H��Q��i��C����Ik����*#"�Ƚ۞3
�mY��	��j��e�o�z� �VE����.b2o�b,��dlo`� ���,?� �1	��;e(�h<��9Ėx��@�&���aRz |�u���rAA�U�	���� �3��k8���S���I�_?�ZN�(H�A�C�~�"�| DU��N�1V�.���S�o�O"�R*�u��;*�M�1c��:0��O>���%�j������۾	�xb �ж���ݩKꊚ�U,-#E�Ƅ����q��ͻ�>qT�24\��(j�yfu�` 9�(�Z<PN�d�����*ɖ��|G�_�J����
���,q* ~�p�R�d,H���~��z�F�\���h!��{ܹfWLP�t��lYc�� O�Ҿ���	˝�]���R_�:��Ɲ"���rG�⁹���mK���2�Kp�g��/R+�d��F�2ZP=El�qТ�a��^�	Ė��K�4׵>�U�nٛ"��w5�|���s4��?F��{H�p�`������3X`�LM��?�&̐?/U�M"��>|�x�D�����??�.�g�����;�x�^�OY3gc��}�j�Rso��B�����w�V����AC��m�C|מ�N.���b�$��J{��A>߯���A�w�z$���:	���O�a�Z�a������]u�V>�/��4��ԡݴ��3U��>)n���_H�M)�<�Q� ~dN;|���ɕ�md?hi�0�����Rr�ПL�Ã��ّqtHn�V�������I�/�}�K%��xL���ҭ��p��}��b�U#J�9T���k`ٕ;�?@����<Q|���ۆ��R���S�2f�64�G���a{��G�~i�� �Rx��i�+C6#�]Lh��a
�}@�Qj�>�u)��V�P������9�2hX6;��*}(��������K�}���φ��+cAC5C��K-�0��6܋�;�S��#d(�I��%�ь�?�nhR���u�.m쉧IqX��>p�6:��yI�n����׮���o8s	q-L�G/�,���)������#^d5T�F��PI �{�8��'�*�#�54N��Ɋ0�`�B��uK8���ej������zԋ�c��Y���O���;'�;M��rA�`d�� ��u>�XB@�A���eob0M?�&[
��'�G_��)�*�k�	�K-�.�ݤ���in&���G�lb�2(���P7*���w
�'Ec5w�sQo���Gy�˲�}��ȕ��;�C=��b�ղ�R���\N8�h�����ٮ����и�_����@�.�p���]�C#�ƾ54���0{����R3oD?���N2�T4c�ɥ�* ?찜+@��;�%���c�d�؅SG��G�i�ٚ8��+|̎���rv��8<��:Z�!b�R?"�j�3n��`��:J����x�A��C)��[;)7 � ���8�S�c��:+� �e]��.�t�Y�]�ur�|6�����s���/ū;H�*,tc�Ԇu�g5g���N�ʉ�E|�U"F=�{�@�+��# ���