XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��V
@��G3�.���ꔠ�st�5��T�ʯ���C/.���g�I@��z�xpW��ƽ*s&ݑ��߫��,v��E{��F�(<���� ^�w��p��YB�W�	�>4d|5������G�l�q�So^BnNO�8��~gJ�d������nF�d��m�km6�����Fx��E���*�h�,!1�_1D⋶w랋�:�ݏh��~ºC6u�OI��+��7�7)��h����[e���]1�"��l�ʏ,�0���RV��;��~9�Æ�\��e�fΐ�͔��i�1�5UF�jxH2ǏX�x��vn?�j�̑�%���.��յ�[]u�G���롍G�-N]ݾsE�OЋ��v���ހ�0D"�4?+8���N�L	�����Gڰ@#6Bm�'bA�k� ������XM�" *(�L�\&��*���YD��l}�߼�QQ�&ד�ڸ�?]J�G���z#cڎ�z��c�%FQ��S����z7D�]�]��v�f��Q��������H
~-���fF<X%bQ�{��Xi֧V�z�cc%���9D��`�g�мb����+{h-�w�8.����O"� ��C�&ɼ_�b�P�i�BD���\';9s׽y�S^��S���(�a4�0	�� �q�v����z�F̘e����H=f/�ٷO��W�Z7�/p+̯Y��dXx0;oC*u�d��ߤdE1����01Ra���7Ye���x��"\�dRk�,�XlxVHYEB    5237    1310[���~9J�i��X�|�$�R�c��Cc`� �]�8���[{���4��T+V_M�`���i�KS����r%I�̞��*i��f����r<�
� ���%�T�G'�b^+=���m�����q�ձ%�K���IO�ۖ݁�.ٓ�r�u���L�T�I�x�YF��d@<=�)�Kة�e��$�W�&L�OL\T-ֈ��i;�vY�U\�UzW�<D퓱��]M��a�n���z���U|%�Ӡ��^�d%\�}��T�VaQ�X�I?M�T<ƒ�=�u�Ջ�W���L�_Uv�XC�|�'�L���
-#����Mk�l*{g���S�_��-X����-��$�����#���9j�R���.��G3��0i�������1i��ͩ9ڜ'��k)��W>�q��L�,3s<�:��*ٵk®�5�,�
�0�p�O,uL�,�4�
�X:���k A]뼭C�ݝe�0�4�+�����E�W���64*X����ݢ��s���p����/����$Ou���5�4��ލW���1`��\� 7�Jld,��S�b�i���f^c�{��D���8��Z�����Q�x���i����v��C�)�P鮪����5���=r�ףh����/m~�6_8f~�i~H�,�לV72��⾡SE�p'�Gt�H�X�-��nf��tz��斉���7�~���ir��)�%%�r@�'�t�b��X�e�� �J'��}�E��ؚ���=�3e�&a�������uW3EP��H�;���>�����������ϭ���q�g�Nq,�.! �	�&�����}t���j=:�]WS#2Jfܾ���2A7���4��A��eB�M L��s��7 ��Z�����b	4 ����h5V�G�s'Z���3�AѸ�{�*"�߮5�J�,�x�kf�/�<C��j}��0�*t>!]a��[G��n�i8��!i������X^�.�%�tc�5��Y$d�U檘]��¥�� �O�SlNE���pn���P�.�$y�k�X�ݿ�CNZ��Y!E��A��r�?�*�H�Nc��1��5��}����M3�-eF���s��e��y�@uu�,j���l6��Xŭ��s�yj[f���j%�!{�������3�7�tbMsVL�u^j��Rw^m�� �Q86R �+D4�6�*�J��T��7�^lv�%�p�Np�}V��A���Y�Sxp�՜��Y��Ȩ&V��B�hiT ��%�,u�զ�R��+�¾�oI���R�����)��U�/�y~%Q>�p����2�&R��ڔ�����#n���cw�"?��ь��i-�M�����	�����F>�=�M�
�(�������" ��M�=������B�2C*B��=��
����"^����,�����a줜&�='�%�ŗ��StQ��t;#)эb]`�	0��}�ݲ�$��tg�Z}+>e��Jjwn	�vlMMb.��|��r7�����qugJ�;��ڗ�y�I��(Y�rA~�E�}��;�wA�n=~�"ٖ-�Dد6G瓁uĚ�v�)|�s�Ĝ�0���k�)��Qr�G�{8]� ��t:��*�1�g�h�{���0RJ\���w>�u���4����权��=�\_yI)�D�!m���-���3~�Vr�拆ΨZ�Y͘�p�h��s���_�C#&�K����sۏ���2�"*���^y��wӑP@���[���(�ZB�DW���]�e�*�J^F������5G+S������w҈���j��',~��X��5neޙ1�!�%���Q\���g�3�/��CG�#�c2D,�Ίb�D�S�_}�B�q���n�4xs!�`�[3C���I�,�y�RZ��V��)��dv��80�z[�V���d}��ͮE�a�%t{�Y�#x21,r�	W��N�6\<�����XS2't[ k����T�vE�+o¡S�C�q���)�+I*��`Q֚��������j)>�谝ۥ���͔�x̀�i+�4���MR�uȧJD��_�c�c���o6<a	iC�\=��	����%��<1c=?p*I�m)U^q���UIS��ф�˨s���a���ƅ����QGΥ�!UU���q�|�[:����C`s��b��k��'���	/M\�j�&q�50��9��&�j�������u�\����
�'�\�	8P��#i���4�\�u%� ��Q�vA'����o����hA�AZ<W�CuI]K�޳��~qE<|x��U�!-g�[¼[XF��Ֆ�	��&�!������6��h__�0�A�L飷�Xx�E�*�+�"�����Q�r�5B?{"�'1��5��{egf���y[+4Q �`h�s�{	�������N�uj����5e}H�s��T�L���a���0�قŭ4>?��d��V����"�^	e�cN����>Oq�2J(�F���?�Z�kv.�LZ����m��~��N.!�3c��'�ņ�J!��UyN,���9��H�2�KW��=�m>��<n�>PZF[Qc�k�w� �� �B����2�M"���i�� �b��DU+��W�H��£̲.�1��3����>_j��G̀귧���tS~dll֊6�F�)	W1��F���h�7j�;Si\Q[]���!���"�͈3�o=�ST�v�m8i��U!9��u�7�xA�N~�kx�d݇�N������N��$���{3H�@c��[��Q�Q���9��^^��oYR(�u��	�.���D�ۼ:ns&��P	�C����g/ļˍ���"? �o�9E�[J6k�}K�y�	�cJ^��h�iĬ%�5�m�w�1�Qi+����͞?�U�
#��*+s�៏ƞ��fh��j89@�Wq,g� k5)�6Ǧ@ڬ�֡��	�z�����уҌ��UF��;�/�Qƌ�ϓҤ�z�b�a�~���X���r�7S�fB��Ut3�Z��,�b�H�w#oB;GE�BW>��D&Ȳ�A���a�貫?l��0ɒ@�)���ו	���g��IF���̞�8A[�w%M�ב|aTE�0r�B�_�3��LQN�0/V�Y��I`���eHn����>�zt��DsP�H�q���4����R�!f�[�9q	��Y�w4Fο΋����Oz*�;�t�ɲ��
73��G��޻JGS�m�A6�(�HU�U{ $�Cɍ��F��$�����-����\$d!�)������	��>�<�iw|�]�����.%��}��w�9�4KS���ű#>��d����x�\7�j�6��Do ^��X:ڐe�|v��\��J�@ν���_���+`u('�����)D5�ߢ8_<(�n�.yz�e��-�|��y���7�i���_�0N#9�]�ֳ*����Y	��[ܾ��7:]�e�*Hp^t����!��XC%1�K
�ٯ?Y��L
{l���ԯ��t=��Yf�e��,�zW1�:����* D�l��+�ً���Tf�I.�0��'x�EH��c����V��G�q�8d}Sτ�m�*��u~����ځ�^�.C��~`ΨZ��s8�:N[�`��|.�%͐�k#�\.�;ނ�n߂��r�x��aQ��cB��<S��pu%𮦾:����)An�2r��S,0i�g��a⻛+x�F�.v���k� R��f�]�"Uϖ�½�>�҂���wm^w�s p?V��~�s��eV��d<����{����\�{�tD����k���"d��͋ʼA͎+������b��"���e����jG���l,��Zz��u�sDM7, Z�(�KV3�7����k�,��J=r���\��dWt�)�s�А�F2 ����
7� �3�}��ru]�㭋n����u<��Q�*[�u�yS?o�Ic�;aަ������9�T����)���~j&�1b0����r$cE��va"�ʳ��0W��`Cg����RߟeX�rk�Z�6��T�KUq�@�;�&��~���K����2Z�Y���|� �%2��T�9?[��b���wnL����ȭPm���
�d��<�x�}>�v��h������b�)Y5�w:�]
����\R^�k�;�p�>�}�gS[y^��8v�xY�&�/�nt����/��qm�,��ﵺ��(�����Y�P��EW�Z��XF�;mR��4�e�Z��\�R��f�f��!���S޼CE�b_���!�Y�[#�/2�@��$p+��G���l$f/R.�y�b�˰��zR�i��hzW�"�VCM(#���d`��ܒض�У%��P�,͊98���	����<��J$oR\�Z뤂���F4!�`j�v
����53�����k?�B���Ԉ ��T�;���M����>r�����$?����Xk�X.�g#5 9�-��Z��\=.;����X��K}�)e$�g�'	)�pC�]�*�Eֹ����zz辊��{s6�;���ݠ,QB�ud�T%�����@{��j~	w3QPh
X�� �.m��!��������)�1����x<9֮�e�����p6�ƠG�"���
_B֐1[^,�>��F��I>�k|Dz1х�WVbi� �γ����+��4Z���P��J��hQz`�x����2AWCi�$V��t\7<����2T�ԓ��ӊ{�ϣ6��ɾ�ڮ�:��xҞ�#ξ��PX�I���!u���Ī8�Y��?w�O�eB�Fx�ݬ2 =�G����0u��-2�%���ǲ��p;�=uh�Y��F����=oF���U��