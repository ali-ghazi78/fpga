XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���ϰ;��ָ&���L�
�cF׹X��nlQ_��u�g�!'��Ž�%X���I�'7u�;1:� ������[�Z�����X��?�p�T?=��@rQ��D0��q��@���U	���-
 _��ȯ�dǶ�l���q������C$��>RR������P=���o����o���2�Y�؝�H�r�au=��Wո�*�]�C�8�t��$\�g'͜^��$� ,D��n���������|"��0�$��a��6i)�pQ�~����&gj��aI"��)�&�"�5�w%$�L2��	����h�Z��n�PٟjZ%��
z����LÏ�á�~��9Z��K�C��A�C'ࡢ"��f���V�X�	OX۸O�&���FA��⬆�aP�9 Ch�BL�R$���I_MԦw�_k\��V�u)���^��Rc�?���c�� �I;��i�4ly1e�,p���ImD��
�k�ׄ�7���o[6\�p�Dt�+���A�C�0�c�:�
枰���w�s�K���5�4�/l��y���v���	���?0�	��
3O8��ӑy��bp�F�MT ��h��ʬՕ�ֱi���>�Wu��s�͠#=�9�}%O4ip�er_�չQ�nj9�����q���t�MXc=�W��)��p{���]E (o(4wVK�q�0��O']> WO�A� *��Dw1��6@xpN��
�vX?کiW������[�IyA�`�"�ղ��XlxVHYEB    2a39     a20�e�f��3�~�/>o}��E� ҫ�*xbA�V���XT���B�so�V��UݸnǽګRF*�Ԍt�A?���J�h��F�!��$���IW��wm�-��V�o5�*�B��is2�U�}g Ȏ����d�Q�ߘ��M�_�h�Ԧ,fQ}iD�	���9�V��Ս� �����Q���#�p1U�ȿum���e�UX�z��M�س��:�-�90θ���Z�4A�FkzB�zB֔�����^J�d(�����F��2�m��q�� WϚal���j�� �b!����7�h��*ѷ����I5I�~����t�
$$�<%�`���:�}i邴�)�(b_�"��S�uw����W	�)ԇ��������@<vGq�V"`bT[tm�k�����+gs M�:d�Ѽ���9u�2[Q�Tw���M��������Yvvߕ������L6�7��Ops:b�����`uD�m���*����n^I�,O4�5}�X%.�,-o���S���_�h7�+Ȭ��9��M�A��jެ�M�M>�	B']Z����A����u[:\֯\��	"��ʊ;Ήk�0rᤅ�]�0��Z�"�L�6M�I��Rg��t�H�RD ׆_W��pJ;
�p]�A�̑��"��P�hoY��x��z�����q�����4U�����Z�K.�z���:��P� ��p��1}�_
x;���p����`�@��Fd|!�N�	�~���;���_��n֗�fWH�4k�"ܾP��˳0\��%H>�t�O�~O؈������0���6�Z
S�e �񺊺������Q㴿���g j�T`wc����N�7�硱*�bWx��|�:��t�c{{�D���XXz�����ʝu����кG��%��H����b@ܔtc�������c��vV^����7>��|���,3�_n��9G�a�K�q�B<'t XO��乎�e�	I�2�rISC��<���+��a٣&���T����[�+Q(��QT޷�c�@���G�+�h��մ��3���F���©���빃'�LT?�&��$���&, *�i_��t��H����	Ce�DsV�(�a\��-�R��60i�G7��dU��Ue-_�V�m
|9Oc��Y_7'+�D#�Q�BۜA��I�U%ӂ�`1�!�T|�<�l�9j���\�v�V45=��
�)�L�{ �9��I�������þ����N��E1�B�I[�b�q��K-��E��ʄ�&����3��T��/���0��I�!�!�����
 \sF����#ʬ�g:0X���(ƕ]e)��A�y�S�Kr�酂�Q�\��� lM�\�3c�A�<�qdi��})=j�fqh&N� �( .Sp����{gx�}(�5�3O�� ��m��N�,�'�`.�'
��:+�s�3��3U���*��ղ360��#/E"��5��ԣ�ޑ�!	_>~0yt�!��%* ��']o��4k�L�V����	E������� �CQzh�L����Sa�:[^���5`}�L�W��������!��fN�����k+��cQ����R���v�t�{������7FLM��/���e�G�.��%�Lᯗ,�L���'��o�Ʉ��1��$�p]�ˠǕ�w�%�GJ�bQ�o��C2B��I�9�o������~�D�u���K�O ��dh�Y^�G�j��@�R��ش���}���R����ʱ�����8���mT����rB	n�)<�� ����브�j����h(
n&6�[�9.���;b/��T����V��ĺ����9���X���|��lW��}�a%�FP�7j��f�<G���9d��hx��h�1��|UOH/�2���T�)�]e�u�����nR����T�����4h1����py5�o��߸PV�C��W�/�e����]W�1os�J���F?�������Ks�X¾��M��6����{�e�7t�d?�������ᯉ%c-
e����MW���Z,���y��p%�F���L���rk��.t���l�%9Sy\��I����I����9��)��A�a�66�{�[�\��cb������,Ί����
��/$�3S�K���"?���ҩ��;Ī1�q����Y�yߛn����{aTB�u���?��*�4:I1�6%��(�x�dd+݊��)'�4��ǔn��u�4��B�Z��Lx	:P�� �1�fp��{�{���gS[�HvOگrm�:.�ZJ]N8�SF��mg�i�d��h<��=�%��W����o'%��ƪ��-F��şҊ�,n;�
�i~�2@�0up�g�=A<}�:��ע}�̡����+%�|���j�����սj˨~��u���ˊ?��߼v�)��ԞGztN��"�S�kP��V�ڐI��,��?ƃ�0�t;���
�����شB��o�#�d�����W�m�� �`�ab^�O*�f̽#��V����'��s�S^����lQo�p�}�@l��TOv���l�!N�i�F���A����[��%��T`���T��|ɥ���!s��U�T5i�;7��2