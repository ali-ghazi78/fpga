XlxV65EB    1f4f     9e0�EҔG}���w��qq�/n�p�H'f�1z�sP;��嵏���JI<�c�5���ȇ@@�I�L���cv����RG����e�\��GHA���;#$I���l�,w:�*u�E.I��6c	�����M�kj��[悔j�5�Y�Kp�6����x�Q�Ύ�4 ��X�W�"�d/����ƻ�2��Vgy�~l>��UA�Q4��'���Fg��T�zAI�}�r�Y[�]�#kUl��߼��T�ܪ,)~���Bj�v ��S�O��U�q����#Z[Ҭ�#�E�ӂ���ME���2_G}@�����?I�p���-��	�5g���!�'��SoC���ni�-�!ϰ�G��a��u������Ꮵ�Ϋ��t�=�|����7xJa�:���Xɱv�D��-�wFV}ϳ�<���QE�+���֫oa���F�Y�ǗK5���PZh}�c�ME��5��maF��WG�.=���\d��/>�h$K����ZtN�_X*�[�Xm�쌵�`�Cn
��̛��ߩ�}�l����dØ��j��i�f0b|� (Ns�-��"t�m�0:˩��zḴ@�Ԇv��Rk�Dz�F��=D��f�o��¬6�=�k��"�RA[ f�A�|",�� c��Ͽ=������d_򉒦:"O=�XP�ވ���>E.����v�ߊ�ޚ�Q6/��<+�Ǚd�:�aE�N��_�AN�W�).��)���y�F��$z?��)���R�p��CMn�J8[�'w�]ŧ�'B�B�ҋ��C��z��U��5d'be�Ϸ�������:!ޅT�T�,��������7��>*V0(Ѐ8���Tx&7���|���B�!z��n��K�cm����'�']x�v�!�P��k�n��W+`6(���+Du�غ����GmuB������d�N�3�n�I�g�}D�%�ǹ�o{>n@�]=�zǬe�G~��t`3A���X`�^�Y�,&��G�O>��F�N�p��R/���Å͵z��|�\9�V�� �	N"gv7`"��r�D?��:9,���g���S3�C}�i�Ć�6n$�,htdR+F�vX����Vض�
˼TJk��iG��vMFA���?�y{+$f���-�L�y$Aֈ�U��q�uU=L=�Rdhw7hJq<z�w���@����NJE,���RNZn��O���"8皃x����q����3�e����C��bo�}�2c���"����	�5�����!��r��ӾN"����դ����[σ"tއ�Ӥ�du0��E ����Զ+MvQ����⡰�;��`�ѢCn�������&���YM���r�{�K^�����"Bi���]�̦"�t�㒔���=��*� �{�f�O�����U�v�-�c�v�2�%����S{�u�v]��Ew9���v��Y��!E��g�$}>g�{@�T~����Y�4[zXi;�w7X�w.92�d��Q��gd��*@��[FJ�K72\�y��Y�;
���-�';��)��/�G|�xx۟�ԶG�%��fP�ySsvZ�V���_{[�������a���]�DI��,P�X��}�w����Ђ�c`M4���]���QʊӪ�@�H]�!&d��I���[��wP#hR�M�J��[��'(��W���7�YGmW�Z���7�-�`�����؏&^��O��8�|�PrR�સ8���r/��5���i`��d��}$�g��h?���,�0���T�L*�a�����_��+�723.C˚��C)&��d���I�[c�Jaw�Z0�c;'Y8lJ������Z����� 'h�a�tg�P�(��oG1��|�qC�@��Y0�A�AS��z���>���4NKT�(ty�<Cq{�+�h���H�\N�ا�d1`�gC�C���C����/l��#vBo	mם*6��4��T�~�J�18���.:jJ�$�[��%�îGZα�O�+ۻ�PQ����uB�����Q�.��6�~�a���u�8B���^������|�w��
V�T�Φ}O_���@B��<o�;�g&��?�{N�����!�g��;��%t���A�* �ܷ�	a��g@.v�Ο����V��������sp_�M,O�>����G]yG�����b?��r�8+A�.*̃:��H�Tbȫ��)))wu��jM��?4�p]��-��e��|���ڌ�3�O?�����<Xtr�Zr0T�����|0+������ 
k8.O`?��v�������[����-m�����`��ŶD+�p4����iv�V��%8������t�]������P�l�Gk��XQK�|�ڍ���X����gx&�?��`}"�I`��Wޓ���+5���ei$yѕ\��>O 7W����
U��Uh횑~(�6@
�5��4x��RT�$
	�_G�Ex�i�{ ���ZgmJ�j��f��8:�rMB��e��K