XlxV65EB    3caf     fd0�s�B�A�"fy�� Y�"J����ŋq��q�o'I#���-�4��x[)z0'JjYd����;���yI֑�H�^���M���'��u�\�b״P���V��JTxCK(?�C�i�w2<2����\_Jx�G���Z�?�ۄ�rj�u`|A���`�=�y'S�X���qx��BYj�=Emt'�f�<C(�	1�n!C����'hh]׎ �<��D!X�:�p���wU��s�T��<� �f��?Q¹��ȋ�p�Ư�ߘ�@��f �]hmЮ3;�>pbeE?1�v��1~h�����V�P�'��#i�
�p+�R���Ot�J��l���1Hd�����"���	���3�����t̤>x�l&��}�uy�'����x���| ���5L��ϊ��8��Ćc�*���9+# ��%n���y���"�[�7ю�����1�\�EU0Gg����=P��ƚ+%jVq
�X����׶�V�<0Ym]c�Mv��HfR����
O���#D3@C�tV7�T��1lQU�Ӥ6,�>�B�DQ7����f��t���U��?����~u��^s{g�I��c]9��۟4�O�k��E�vX8�������.VXe��Zt�̔V*����
��cr��=��)R�ӿCu�L�у�6G��nm�Z<�=^����8Z�p�/>:�H���(���5�9aS�(�/�r}HoҚ����X��s��,�k,� ��sM�X�1e�R�r�ԞE ,��>9����I}�Oڄ��K������п~t�l��I�Z�^4���\��#���<7�5x'%C.\1J_��I��6���v��L~����B�����I3���j�;R�ƭM��ÒS��DS�4ooc�!��_ �yֹ�5�F1?�������W�A�Z"���[ !�G-��|�p�0h�Ԏ~+on>[��XN�"���p���(�O�;ّw��q�-��u���L=�R�I�'��*:�	o5�{z�n�Q�d«hWF�^�)�pѤ�k����2I��\Xț�hV������";�ߦЫ����YƗ��H,�+=�B�ﾨȘ���
�{�� E�hX�����Uu)�}<ʂJ���$���P����$�5��֚�k�r�����H˓���ޙ�$o���R*\���c����B$�,o��}/�t.:�b�����I"V�զ����{s���W}c����������DX�מ��I8��\U>%�g�pZ�~�N���K�����A/��a�n.	�B�д�谦[�S� F��W��ns�t��Z4O!���~$�^�E��88�)Z��Yn�R��@7� �_��ÄV˪]�9G;�h�@��Н���3
���:-g0��ek�B9�M`گ�8Yd��	�%�/s�|�k��@���xx�(���6f�nk��}��{�
�}���MJZ�jFQ�������lG���ј�T�Fɑ���MHK�3B�c�QWR�����"��� o>��v�74 Y[�x�k�|��v���uNxݏؙL��
�5��(gg��D�|�BC��~Ԥ�(c�Ōx�	߫�cΞ
@\�HO�1�^�0���ʓ�1�ߛ�^Q��H~�p�{��T?��Qa��Z-8�ow�B��ԥ�.*&�p� �r ���Y�(s�����=������_u������ &㲐6n���������/v��i���wS��[�ʻw􍪢�#��٥��HVh�|8�FhV�	�a��j�������4n&WW(8�˞)��!�٠'����BT��9���S������K�T�y\�i�,Lǹ�r#Q�7m���"�k��2��'��Ђ����ѓK_���O�T�,���3�r�t�%���u���ad)Oo�R'�����N�\�ș��Q-�
C�q}�-����T��Fi�jbp�h*�ѡ�Y���A�:���g���j�avXZc#�WM�Mlf	Ht�d+����Z��X����S�k�.>��R��؍$��n{*U��F8yJF�%�[���P�12�/PZ���&�{S�I�Vѳ¯��i��uv]��@$�P�e�M��z�հ*��>�|�	�o#�t�\�|B��c��X'�N�?qw��0:E0� �8����i~8n<v�O ߳f�_�C*a�|�����\�A��Qu[��Lִ>�iH�#�P�KģEơ��S�hc�.�=�� ��ә��1�y�l�����Z:�}N#G��BU5t�S.o��-�p���*�pgFB.�i9�i�g�������;�2�F�!F 4��;�V'����@JU�b�P��l�<<T��Z���&���[�I.�QZ�ّ��apO�H)�t]`�p���k#�z ��B�c�A�,���X�
�w���~��wՆ{����y&���3��7�p��~��?����F4��^�m&v���<�1��� �!�\�he�sRF\i񺾢�7IǮ_"������N�l���`�ar�!t�e�ˈ���S7�p��`�:T�w�y%,�m�����o��-)���x�{o�ģ��V���{+Ȭ��Xzx�i4�z:"�(�{/;�������۲�ɑ;j�H�����c!ɟ;w�N_�9?y6eq��%vX�ӱNv��N�r{��U*�b԰�@��nN����`"�Ӻ�N�#�l��_���xU�|�Ne@^��.���{�2�e��^�+B� ��D�NN]�F��8�yYl~����!4���yq�z��sƒ"*�rrd�[A�(k%���X��er��3@��/���a���>�1=;Sw��:���������1��yeZ�Z��{cĵ�me&[�D{P���%�R7n�QL�(��(V��;=+���M`��9���XE�d��gPq5c?��� ���>Q��n�����T|xM��+E�Fۄ��>����N;ͱ�2	����֭8�� �u����4Y' ʊ���:��K�XV�4�!ξ��a5�`�P��`Nh���+kAI�f��f{N`b��z�!�SD(�^֡~d�٘��G´�T;�$ }�O�&�d¥ܢ� ���N����@>�'�s�ai�|�(Vz���+�\D/���o�R�}Ei�������lFNk�VL5fW�5 ��-�u�1�O���8m�`O���q�s���|�VT�ߴ�2�g��G��l������%��S��NF�3e�=q������_�V�e��дN��P�p��D�l6-�:�Z�)��t�A������ȊHS���ad7$���Nt����A��c����q��('k�[:�BB��fd�Ke�	T�=>�l�7fǾ���4���]������z��5�<��*����3���C��%%P�e������n��氾(a��O :��dms��bQ�K��W�~��e7��L�mH�Ö��1l��U<f�N�AU0)����D2�9F�UUKҋ�V�#�I:�x��h��2睚��x~��n[nL;X�n#�%��b�a��B�8�����~=�&a;�(�٫Vg�$U�ژ�娳�6j�YC�D O�i�I��Ӹ�0�D(n�86wV ��3�WY5�؄>���HR�^�][L���ìq��j�5�ofnK/���ͬ��F*S��7WȽ`���G�k愐���R�I��:\mo)iɛ�]>�������=�}H���s< ¾���9���N�%�'=J�q�,h��`�T����ܻ͞h{N����xj%��]?6��]�R/Z;b����-���ͤ�E-�."�|�a��Oh��[���=�=��G���ɼ����E���#�2,�X|>��iR�n����t�h��@�a@k��i�cS-�C۶�	���JHt�Mz�RO��3R:a�<�	].��=�*�m����� R'���;nI�K�UU�6�d��������v�o���ч�Q���5C���@|���ႰD=Ї\�$Ѧ�a�)F�k�ROs���3