XlxV65EB     81c     270��YĞC�u�Q��f�s"r��+8�� �x��蓹N��s�l��X<���2n`<������.m'D ؿ�/��n�XtjX�I/	��Wv3�+�C�et4G�Z�v�XJ:��9<��Gev�e�,1���KI�WP��W`Ѿ�D��}�D���	�����%{A.'��[z�~@;A`8V�k���ٗ~2w��T�`=�3�e���&��0�Ds�sm���`i�DLj0���Fm"��f�S۰芦x�|�D����+b�*H�μ�fy���)��#�b�_EM<`��ǿC\pͯ���j��3<`'0|k)e��-�����f,�8'�;����X�_A@�jEqm���Xq�	̝��Y����i��Տ�fH� 	�>Y����g�y��[��zs��6�&j{Қ<d�I��QE��ů��C���"�u�%�i�h��%��w�^��;�8VſV\� ��`{��;���&R��şC#���|@SG�c�J���7F�\�3Hf��8�\���IJV?�T`ʪ�������B�ݺU��@䃒{u�֤іx�R���|���ӓS-�=s6Yv%�J��M�; h��>�_�LȵJ����1�ٴ����`Sl�!�e