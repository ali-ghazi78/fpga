XlxV65EB    5145    11c0U����*8���S7QD<C&�̧��RW���Ϟ.� �i�U��R�Ӄ�ޥ�+�;��P�w�m9cP��"Lg���L|w�̵�D�E��E��;���J7]����OdM� 4!6���G�x�݉Y}%Wj��U�$�䱨�L~M%� �ˢx�� K '��zWr2�#�@&�G��ǰGx,JJ��?�~QC���ۅ�1�Ue��/�ea?�g�W� SȀ�����m��oXc$�E�2��َ	-B6���ʃ_G2RD*a�6͙N��^''S���p��@w�zlłx%b��v��L:��G�4���R� �5/l+���
>U��9Ŀ�<�tC�K �vF+�xE�L����]CyP�8�B�K�5x�G��	�S]A�;=iw��s|C�x��m��#�$6;{ru2�}e&񍂸Cq����6�����2m`=��Y�Oa@���T��
�٤w���|���f"�A<O�X>]Ӗތ�Mg�kx5���_S�� j�Hޗ�k�G���`H~=i��&��F=���~{���5��Sk���[NJ+��gfg� ��=g�:������"���[��zb&@��})�ͱG�����4�%ѧX$�3��P�����H����xy	/hNWu��=x� ��%j���`2F@��J5��-�gR�qȶ�tN���r����צ̬����	��r�0�P�[#N[�Jw�\�Z��8I��C�&}���"�-����q�|Gg��1�\\t5sHQ�����ɍ���Sꗞ�Z��bg�;3��B#�+������d?}���7�~���m���JU��N�à�N{����u�"�Ov��B{R�� B�x��zG�l�U�`ٿ���í� ��6�@�@�L$6qr�O,��E�MW���3�)	�4��)G.V��+�]ldE�L,@vd�L	k�K�d�RV���0��0�� ��Mۥ��a
 :�a��sP����X�ү�~S�d1����D�\�tؒ��jB���O^���� 0�r���=2�!*KF��^�A"���'��ϵ�
�+�����F0��;�����*�O/&,儧^�T(��d���˰F��b�`��QA�]s]z��yȀ�]�$	�m��;�<�M��9���{�ռ����*��}#p�,��'���D��.M��5�����B�Ja�"�s��%�W�?')�C�{��%5&�� �Ȱ���P��'�U�0Oa&g�w��j����q.v���SG�Ő>=�֡q?wLA�tQ�8�1Z�W����I�p~�w>N5Y��
�w�� ��WA��ڬ�j���?u�Y��AԖ,z�RՋ����D�w?��ZʭU6��j�4r��T���יx?��1<�`�T������sx�Z��T���M���ے��m�i,	�|�F�ql�lZ��>䜘po)����>�ѵ�a$�K�/��\��G�P]k }\�_�������۪��(5����/��`Ebg���h�yG�T'X���14�?�v�eIm�&i�jB9.9�A�Jz�7o�Q:%'�� ׅ����"M���,�/U��{�G�`ٸ�|��a�{Jq����t)���t�ZH�����i�x�!q�D��E�����VFka	�A�\�3>��<�>?<�����w����^�8��7��T�
g�6 8�z�_����o�S��	�ߵ��M(�4�:���{Z�09�$��n$M�{��;|��G�
���zx�*Rma*��mt�k�1�bTN�N�[f�0�o[�d��s�k���;��G:������rN��v��ҒQr,����Y�K��q�p�Iov!�Z�QhvV�n`_^��^Ӛ��@��Ԕ[>�r���ڪ�!�&�J��?�.�M?B��������k~��u�=n���% ʩ� H^��D�1$g�W��c�Wjy%԰���Y�4��ֿ�פ��䌼R>�N\�I�@�b�x���}1�Ö�L��̐�/��iN�/� �g/�#d�߶�L}���[VY�f�fi>�6�� ��S)�Q��ی'��8��4����ʐ�
�O�̆�v����+��l��c.��0Xl�s?,h�3�|��b�;~�4S�ޘ��+MВP?k���+O�6޾K�!$��������h}��[h[!�z ^��*��C�9������QM"�YCm�b�!���M��
m<I�����C��MW�b�}�E��GdY���g'�G��Y,�ʢ9H �x_���˒�H&T��:-I[�0�ZHJ���^��=_�P6@8��vd�2��~{�W��m5�&��<
���j�ܹ�)�
���-9��*O�knt���O$�BY�`�a���:����׃�c-�`��uG%�!�vtL����v:]�
���G�<jE�8�A͎Lx���k�"q��_z�ur��f�a���8q��m�*f(o
�!8�' ~�`l>����'Q�5�[p.6��~g���9s"�zS ��^�ͣJ e��ו]hVpA8�Q46=1}m�<{x�A�[ ��J{�ͷA��:uSu��_2]�gh����$���7���A��z8�l���V����~rꩋ�&m�#�-������{��"�&���S'I��K�>�ۻm���AD�Ւ~ ���q��b�% x��ດo�5X�l������w^�+8��b��� �@K����k�b�Gt�ޮ���B���g~}5�0 �6��j��v��U�:�O�f$��S��\%�����h;x/r��o3���c�ʡ
�J@�F�N}��C"M���A�zm��0�} 8�Y���c?��b�;��	I��e�[hR�%��tu�{��:��e7�ʙl��n`�.M���;���
@�����Նjiڰ"��)R�� �5 _C�ӗ�%dT��~���%�W�ʋ��FY��$�]C.�k1��
&(F�\�We>:�0�(�Œj�z�/d*P���݆sH��4<�=h v��2b��s�u>�D��ӿ~��W��t���!��EW��d%hC���p�jo�����)� ��[����wt���R��e\������v���0K��Mq�ͻ��L�\N��V�Mٳ�#$D@���mq�"R��r�c}�� ��!��ӑ�$k���̍{�
UY��|�4��������. !:�qъ����錇�,d��5W�"5��E\��U�->�����_�T�.>G��k���GNh�9�V�Y^���N,N�b����j%(�'�(��;�\P�����2��'\���&����W�s�)��D��V��ޫv� �S�{S�f�ϛ��E��Ŵ��rU9�oI��zzX+<F,�T �'9 d�eT�;�#���[�Ѻ�US~I�z��J���93�^�D�j�u�wH�fS"��Eʸ��2���t����̇ Н�6{>�S{x�g��_ە�1����-1�X3��!�s�`^��$�;3�t����[A�8,``�umJ}Z�߽*-�\а��F�	,������Ti*|�v��ri+���v�+�&�
%E��P�l*W���7:���U���K^W<q��?��2�C�R�>����o��V��3V����=J�N����ݐթY�����o���!7͹VE�顀�����Ƿq�����I��Kܟi2���G�G�	�ʔu`�J��K�u��v�I�I�f�DE�l�S��t&+�E����-�OY�|҂m>�f$?e8�4��Jc��l�j��@o��?&-_~��d�tc�v�q}G��N�$T@U��b�&���;΍	|�h訦�0狘��;��P���&F#ߣ�u�0�Z5l~K���Q{��z��u;��z�������~t(��y5�(z�A�ٳ�D�P�ܼ�Kg���`�޺��]�m��/+Q��>��0�aպ�CcT��d�.&�$1,�[�'�[�go5�^q�;T�cv.�����%�E�������+~�p�@��$�&�����^�
����G��ਪ��3���\�N=;�Z��>�2-��̪Qݨb�%�f�@�Rc �e# ��
q�=�mA��m2�9my���9Ġ��ቓFd�z
o}'ڔ7d�ʀL���Sd*�s4�G�vֺ7u0�s���6�_�ߪPp7x@ 0�2�Xa��O��yx"���\�aR�si�O9CP��*"X�ܹ�;e�۱V�?�˶؆9 z����9*�|iX���_ާ�-ڍ�Cv�,���9�gƇ-�ۗ��������#�XUm�A��d[�����Jm"$�0�3�?B3o�������L��?�(��q�J��_pΖ�G�6u���]p�GS�d�9"fT�?`�x@���b�ң�h�J��7:N�f�u������K0v�\�g�m�A$��)��(�Ӂͪ�@��J.���b��tT�K#�����-m�ר�q.�},)�a��Y>�����;R����