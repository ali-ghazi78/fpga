XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��@���s}j���osG��JޣC�|�6�/h�}B��8�v��I��`c!8qz�)��پ"5��/�g159�1��1+�2��լ*fҽ#��6Z�#��P_�tm�����TZI,�T���ʾ�Ay;J��|�L����P~���E�tꦅ��P(���3V���� ��A��1��[(ͅ�!�x���f��mJ�
���[��,ݱ�]#�ؾ�^��	<#[0�)�篻�w�>� ,G��D3nt��yH*_�g����%{���_��5k��
�/��`0�O��7&��bY�0�|�?�G<���̆�}JD��I'���H�K6�T��S��a	�Sf�Z��;O9̺��Ϯ�g����2 �<v��Qč�-�e�v8N�E�J8sT���B�X��Ǖ�r���.vFƕ��y�V��B��ń��h];P<�I�58UD��i�0�]� 1��H�e�e���'��sL��{{�����if����Ǒ�jw�|'������`����?ƍ�!�eB�;h�7��� jM��fLRR������Lհ��J3��B�)���-bԪ��ڧ�9> ����	���B�;O��:��S��.6Ϡi
5c}�q�a�b�}0�xϷ��0�Q3��4L<u�)dse~�c5�N�Xfʝ�m$n�6�����}��ɰ��� �������c'��;&w���d�J�%YdG,.�4��_�_�] ��샸k�%~|aU�'1���5n��c&D��1)[XlxVHYEB    1a29     960�����}Ъ� P3�ijxο�",�E�wwx�v�=�������	jF5���!����x9�
7)f�؄(V�sÀ;'Hă�z�E!��x�����C���H#��h��tQ"��VKTq�;5�J�ൣ������(�:@������R�P�A��6�����[MeW��y�n0��4D�LLK��T�$�:�����3��e����x�q�cauJ�,�W~]Ǣ2͚��L��G�&��[���T���������z`r�͗S/�ι>��[��|��q�:R��:D�-\��A	%���*~7�uk�����<����d�nO�[�8���`C������ZGv{?��{� @�'�ʲ��TM���x���G���j`���-i^%�
��hM�<7��U8�zh�e�v�A��4�s��}ޢ���_�>�Dn�8t��~U�$t�(��?0t(��ĺ�h-ʞ����NT�ٖ�lꝚbzp�Q����H�=\Ue,|�p
��O�& ]LԵ�%*Dq�U�h3�jo����g�2��k!�����o�IYG�a�Y���aÿEh}���ިJw�FL�B���K2����c���N-�5Cu{�"��\dp��A��7:tZ��{̸v��5F�)U����ⷦ�p����t'�C﹅m�4F����Z��b2�嬇����'������#�t�Tډj�azS�@��;��u��������GG?DO�(��gw���@QX�:
�U�ky�a�*߰_� Хu����O	7��J����~|���{eJ*S⤘�8��n���H(r��`�[��P�Y��������D�+�}� N*�:;�,�
�Ė�1���TD�0�6JH��a�c5y�I���#�U闄�h(Ӫ[	��kI�!2VjL��vY�(��M�ԫ�#�=�Η=��Bm"}��rf��lV`�QQ����0� ��	ͅ(C�І�Kg(wɞ0��6	"���'-1�9�����A��Y���I��.��T���g`�&�;dY����^�U�ӳ���]!�
K����Nѹ��@���˂^��^�Aߍ�¢;�vj�%��.��}�x�̇Y
W��Y�
�YD� ���0�(7~hS�H��F����O����58�Q�pg�R� fz )Rg ܾ��BC���A�>�og��->�
(��.?
w8eɧ�c$���=�8*,[��Ϻ,�T��;1��Q�ɔ�S�\��4���:�&�ɼǡp4��A�L>�y���?��;{Ƭ�*�6��1F��i�/X�"1T�
�����cF��9_b�G���dL�&���K(_rT�Os��/�0&q'�
�}F�!p�7��sL�!�p���*���)[�%s���|�����9���"�Oqx��w�C_���9,��+\�M����t�=r�@���IjX�o���hs*�wy0)zU��@���'5��[��*ꉠ�Dur��8�C�p�e���w8��y[�'|����-��E7��v�mr}~���blxJ�P�8}<wN������0��;�oz��E�cS`r���9���@O�/�E��ɳ[6��aA���Q ����wq������bZh���� �'N٠�R%���[�{���ȁʞ��|�Z乿.߇���3q�"�l�y�?�����W����N����b=�y�0E�`m�4�y��6�\$6�P�Hؙ������'�}�g�}�S�<,�T�L�Ϥ��~��#�=d��X	�tG���]@b���7~�k�R��X�I����uA
�kz��k=i����u��Td�����Q�/��G�5�()FT��5jb2eΑ9X2p��H:�pb@����V�6Tkʟ�ɮq�)�C���!k���ߌ{`?��Sg*>1	�9(��n�O�O��?}gL#F0<h#!����=o�%��4�m�L5�`0|$�B���w��� L��J<j'{�g��|q�+���Ô��`��� ��QU���� h�8�݃S�|z]�B�p���IkPn��jUS�U�>{"�G<o�1�o���V)o���gi����zv�̟�=�'�8q�͉I�@�G̽$���z7L0����kJ�I2���@ O�����͛�j�Vߞ~L=��/J�\�oᩖ�ĶB�;�++�����W��ŉ���_T�ztv'|�l`����ن?ͥ�t>N�Gl�Y���Ttw;"گ2�xʑfV�Ӝ�A�B��R�J�]IzqA���E+V���2A�t���n�M/{%ʌ�)���K����G�ugj�?�\��1��,����/�䖚gǳ��|�������