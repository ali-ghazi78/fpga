XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���vIGy<����Õ�;��QConI����D�;�)�x��Π˽6��bS��V����@�K#�#���g3�5�277��T=M
�R��4#'�u�̓F��{N��(�H�S��U�֌"�m�!�A� ,��v��9�tE���ت4FZ���5�z#p�*y�)����k�����ɮ�|�Ȳ�F�m�8�md`�)82��_��R���
����*Ae�x��Ҧ����=�@?��vME�ͨ��bq称w�R���1BC>��n��I1ة�sP�[Efn�(�*w�S�������y���.�˷�5u�ډ�sJ����x'�L�	��{�� �p�T�ȶ�(6�*�i�R�8b{��)��oZA'ˀ'�CD]97^�ٯb7�d�c�����bL��(Mt�����J�����]��M��74SEmv�K�8tbO�Y�t7	Ge%J�>d3�w�P���
�c����WQ�Uy����# �����5�����I+���F�yU����pq���'�3�8��/�/oR&O/�����gyL��m�����} �+=�j<����`<w����-2��w��v�]q�{IL�W�J���܈JGTݲq�HVTA�]�;(2��k��ӡί�c��L
XFRβ��-�>��]�Q�JmG�R������U讖����;О�E�w�K^utO���v���j�^�@ֹ��'�_�u�h�_�]��{�p��d��w!tyq �Rj3H>�81�Cӧ�~�RN��XlxVHYEB    5146    11c0�|U ���!w�P+p�Q�)��?���$2�/�����.���yLb1|�~���ξ[��j�9�<	ݛ<�}_��r�WH+�5�#�k�<y���"��bY}n�AV��ݴ��FD&�'֕�i�"�ۗ�f�C�IH"��;y��6�DLf<��,�2�OO+R�;�3�~A  ��?<9���3x��
���DAL���r��Ʌ�4�jxk(3\�7?���v��V�鍡Dw�LK��9��-*b� .�;��Wx�F� w(��D��B��Z��rsf���׍����+�b�ꄿ^�"�R79|,���}.�f!��iͣҖ�so������ĎA���vs>�����}���#�<�#��	������J}���֬�A���P�I�J3c�����@{`��d������L���VB^��lǹ	�?��&K�,�����#��#�^y�;e�{���YT���*n`��l�*b7�I���CM��+ @R�_��)1�_k�t��0�4zL�5�a)lbE�`�o-��O�u�	�i�߼�l�����r\���	�9g˨�iU\º�<�
ʭzT���.��g�g/�ƽ����A4�~�IZ��v��T�c����@�.]h�7�B�������	Y��sy��Z�dE�Y�.j��oRnj�j#���R�f� �����k�����Na�~���= A�>�)�Z�@�zD��F��a#���0�QK�w1'[�P����a�@z�B�܃�Ӣ�%�
�e �G�C�0��[+^���� s�R�}�0����-�/ҶV8��&Mq��4��3y��I���C�u^MY�O��}�����;x�hh���ygr�t��r����Z�"F~l����H�R��z�AM e�/��	J��	4aO.�zRO�:-�}��5�Yx�8꣎ŏ�F�3ۻ�r��r(�q���ո�aR�ZL���mؗ���Rب���P��a���(��I���L#�:�71o���t6i��o��� ��B]�3�
k(�ҍ�I\F S��5�n��d^9�sE�2��΢�%����G$��
Q5zG)C"
���,Yh��0�f��q��*���;�i��������ɄI
GmS�|�@�X �c��R�qy�H��
�5���a�d�s��-�����Y�PL-Xy�p&�8[\$��ӵY߅�qhcq;�a��}���JԤED��\�$���i��u	�B6�o#��Rõ���ʌ'�m��0SP�M[�z0�uɉ���&�#?��a��}`{�Dyw�gn���L�;��;��$6�,Dio�xmT�X�� ���e�������8�to ����������-���зi�Ә��O�j�J7W��?�`����+HZ�R�Ǿ�0���5h�~9�.�H�x�$��УL0Y]ڹ!��,� �c�t���t-��k�H���Of����)0���["���Ey�>�K�葴X�'<��� �����&�͊��/�Â>�r{���E�W>d^$��&;�I�����QB����;ym/�W�S�b!��4�;�Թ�sEt��6u����;�z��[#�;�8b��`E?r��T��u/�g4s,��EY%%Z��q�k�Ě5���K����Vi������m}L�E��L\�-6�bj�5
9^����RK�w//4�":�d�W��������N� �ԫ+Pq�^��<f���:�"��
�0Ş:)fO_�6u�~�4��zEi�.`XU���|r�FD�u�|C.��k�����L񰳚���,�\u��+)�t:)��6�o���I���8�IE�9��=据���j���рֵx]i8P���#���
T�N�GT��A�"V�]�y�d�����\d`�F)ΚO�C�{��}��^uUS+��噰�T�un�V> ���!���Zm�z��c�M�����*����֜�۱pf]�VsL )��rO��?�nlۨ�:���&�����9:��G�\l�:#;�u��f&���@B]���D"����De�Z:Q�ͺ?��J�u����p�C��/�,L(K�%pbD�����r#O�n%nE�c�Ζ+J˝�i�tPAq[�@]@ HO���L����c*� aK��Ů�0Y�}d���=��{K��;t�����b��e:����P�MQ��.=��۽��.�A�kn
���,|�r�z �ʶ^|x�4�Qד#|����q]��ɮ|���Iժ��h|��W�~�%S	��0S������h�ĸ�e�����ɀ� $+3e~"�biFhK+�t]2��V���(���ӎ���c��zM���.1���$��M�"�8%���Bh_4��
��^dK����{�԰5n=�����&�(Cʉ�ޒ�x�y�ʘ;���V����ru��k�P��0Y��M��w��J3��SC��H�=<�o�-�M�#1������-(6�]w-���p��پ�^�)�0G|�t�v�\[��2S1�y30Z��������>�dL0�pg�.+�	R����`�R���OT��? ��{��Q�goT	I��m=�}  Ib�	*�|�A�� ���� ho�<��6�/�q"X@K��Ay�%��_���\�~���^���M|��t�v��Sy����b��������r�N�Q��κ�Rc.m��CE�]F1�z�+.��@Wɗ�ɋ�����ENbC�F�SƝ��5�[�T����:Z��)�k��8�V���2v�w��at^��e�zs?���C�4w�|��7@1��KA�?�T��H���}�b���D4*�46.d����':P���X�ӿ�нIh�b!g+�e�s^!
nN��h�P*�4��Q})D.dt�L-[���L�����msq�2�aj�ו�PAL��%͙K�2h�43}W��vN5� �fY��ǐd܋z�Ms���â�.�?�6="���Ə�W�D����tL��%���U�f�e�<&����[Ox�ت��D7;��mp乛.	�}���[�<I��"�3"�d?)�ȴ�"��̼/��jh��QH��V��7���:-��� r���c|����T��{�S߉�ߪ�Yo�0��X��<�~q%�SȞ�3k}u���YF�rK�Ǔm�տ��ۍ0������w��W !��܆e�
 �̍��]®�`]v��Dx
��n=��+~��/�frK�7�WA�+���˴Ud���8,ǭs�m�s� <\3Pꌣ��(�J�H�:Q�b��'�M@0zÒb��I<�jD���UX<�]I1߶.��r�2d]��"��8����jvh�t*�u-|��,��g�D�n��ܮ�F�^��	�錖h�?�\`��,�A��`��;�^�%���Q*M��J��*:���H��❪]_���e���� e{ueq�CBy��E�B
����v:�B ��iX6�1�]�J�Ug)z�7ݶc�j!	6��%f�ǂ�3	FG����3����H��h�I������[����M&�\���&�։���y�v8�װa�q�2V�=?�O�I^�+~��,���&�!��9t�c�����E:4�Jm��!�����qD-�.�,l ۆDf~��Z����2A�%To<Wd���^~�/9�E_xi����Y����f�ʩ�4w��������-�ף����ы@I�r��TN��6���dW!pwW��Յ��R��˙u.6��tH�/�� ��
=�`���zBI��4���CJC��)ÿ�"�v���ޙ?�K��-I2���?��Σa�쉄�"'䏡��ؿ�ªoؔ�m��3a��ƕ��@{<)p�P�����@z��"R����t)VL���ec5���U����7 �_����w��)FJ[!��s@��K.�-*=�Jc�Ad���~����+��d�P��̵�7{hy��G9lyyS'�	�������<�,�02H��1[�c�Z��L�l9"M�R��}%'w��U�c�IF+�%	|��xIYN�:C�ٺ��!�}S�=�uV�D�XE����Q1ٸ�O���&������͗i�d��;Z�ժ���g˓\�whU�b|QY"?E��&���Zv�ʀO��^�r���-���v�W�Z�dx�E8W�R�	0ڂ��I����ĭ0eϴq=Zĉ}gwV�S��7Wo��֞@VF��g��Xǜ�r�D������RkT/�:V�oI����m��	��[����3�D6Y>f6�3��3`���N�|�.�{ڰ��1���O��3b��%�LMS$64�؜P
��M
=A>)0~H-&�oF	$e@�=1�r�]�,ÛU*j�8)z� �����z��叇�ʛ(Odw��0t�m' 4D؝��s� �����K~N��]���(G�`	�+��`1���|_GH��^C
^�oq�D-��