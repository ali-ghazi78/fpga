XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���>s=c��>��%TĻ���cL�?!�%)����>��P�<G�| O�<�[�]DEC�������} �f���u���%�d��(/���o�HV5Yx<`��|F��`�2՛j��+@˫�vi&��h@5� ��6�06ix:icp*p�jsC ��c��Gq�M��� q���]E�7q ��:S�e
�^oFM9*��	a��5���s�ꨡ�@@̲F�hOV>D���Y�;��l��:�����L߯�v�!�	;���d�����`g�ߓ�]6�a�>yM���	(���-��a����}�1�W�F|���]�� f�����'�wTY��!k�WH5�猪���������#6����e5�ղ7y IE�ߔp�פ�߆[��M�w����T��6����e�X9�1�7\��{�0�{n~i���3�L\�����r��&�i� �Jx��@�4՘V��͑Fz���SI�i����G�]N.�#��(� �3�Nߞ�c�[�Zzol�퓁�Ea���`��ԛ��QX���3�tKu7z���?��O����<I��V</:���MZ2%�GV�d�#Oy��p��E=E3��,nɑ$
�ա����uBb؉��Q�Ǹk��������C�J���p�-�>!ޅ���[��'8J�@��Du����1�$��{��\����۸�o��Q���!�Ul7�J�d����AZ92�/{���ǇKi/	�F>��7t�qA9�hy�%�XlxVHYEB    3cb0     fd0�2H�M?q�a��k߰����x.r���W�e�-"������Y\���+KL] ���H���
�I/�5��듢�`��J��"{P�?ҷ䩉�͒��lh�4 'A�y�Hk:6��|S}ts�ŋ)���_�91�+��TZ6�9�_�Z]78�4�� ��:0hE1�[�5q:qf�3�?�]�r�2 ����l^U)T��QQn%Q�~���_�����YD�z$���ԍ�r���&�d,���GԊN)hu��S8?e���C ��E�c�^(Y^|��o�p��_��=?8���+@ݴ^E��neX�p��t�xa3r$$+O��>���N�H�赅� �1O���za�Hj��}�]����9`�ݷmT>�*��,`�3H)Ť�
��:�`������=}���Gd�BHz�����G?���7���/�{CÂƥ�+�MO��\ ,Ӯ��)(�1���t�䞚w!Ѽ����eV^�%O�!�H����>�0�q�Qq9��cay�tl�-9Ŕb��IGUZ�5�d��Sĭׯ���X^����3���6�H���p��7��3s�� G�Md.��}��F~}�a���u�Of�֕�
eA�Ȗ�ј\!Q�� ]V�yU��HU�o��eq�5������<*U��;��6.By�	$�$d�ff���`<�p3#i|��*�Mt��.��oP�x�Dص��Y�^Ry�#���J��+�e�!���g�/�H�ؕr(Q� z<i�	��u6�����7{�>s
?!�H% ��LR�:�k����F��<�r@�0��[ h�j���vȢ.v��]5��X�(WO\<��L�H���ε}�1�8_���W��6�.��5%:!��ܤ`���3��Tv�W$(�y��!9��>��0�����U�A��ￎ�s}1��lw����ٵ�r6g�R�w�����\�p��Uy*N�m�
񓃺m�� AfNU�[�>�㬁Đ��T���t��fӂ����m�+eu���B�|�a�[6��
_��\T��I��^���I�W� �I�i� ��W�}�Gj��#B�H�����
�׼��4���5��1����ko��A��pNq�_��io� �T�pj�Q��f��e`�苸�Q�UAc�ބ�k�@�iӫ6�h�m+��PF���fAN��I"��m�A7�h�G^<���kra�����V	m�R�u��|8���������F�?�x�����O���y���aK��|
�����&�
�K�o��hg��$����0u�]�.�?W�1�)�w���Dhι'X��f-t1�2����0�l[ȱ`��9�׀Xj9z� �T4^�Z�%0MN�p(�Յ�hN�ồ�6-%�u���%x*=����^�Q�e��R��ٰׅ���z��\����#3D��of��W8�$�Ow,�B�v �����#L����;�������J���ֈ�
DPp*;��,7Y��kBAr9r��g�U?��~�'<^R>�Ie�p4G+"p�#h�}���Pf�9Ht�1+����Z�Y�|����ּ�c�'�ނ��/7�v��t��Z�!�!5d�Y�����}֋�(p2��l��&hN0f�� ��

į�X��пH^����(R���Д��$�4��V4U��K� ��8Ӛ-@dzj��c� ԨB�]+�M���H1�͝��:���Ҩ�
p��~pE
���fHȍ,?��4{��P���k8J�H
?Nd.�u,.N��v��j��
~��D{�>Q
$5��r�Pv��Z��+|:��57��p�� �'}�{\�K�~ЏF���䌿���s�f��gD���A]�8�o������	�P*bNE�d��T"iv����S\��Rt����}���鵒�h��L '�y�ß�P��y��[�����(��V�5��Cd���8�/��e(I��G�j5}���~�����{�k�I�tl/��#��T�ޕL��4p��o�J`S/S2��W��� L�/`Vt�owC~��V�����k�G���\� (��;����ت��Ռ�Bĺ�H)e��J��H��}i����}��m�ڍ}�6�T�?��u׹�~��_�bg9����JF)\�v��B-���P�G�;�[hL��e��4�B��Ƚ�@#E��u�f�����=�<��/_ ��܊�gV�`o,�j��T!�Ip��E�Q�+�TA�GI'�gp�<��=D��E�f,�\�ݳ\Nޛ�����P��N���U\�>d����"�?�a^�!̘Kp ���h���ϔW��PE�w��	�)W�j>a���G��8Ұ���[��� F�O�����7;��3po��;�qj���E�^��;����C`:'C�����u�x+Jj�	~;p@&b���,m��	/�x�?[V��=2T!1�/ʺ��i�C���GZ�5s�(R���ŏL�8��ޟ3	^Å�pϹ��A��AA�_zR��8L=_m_|;�W�?Q1�!�¥y�t���/#�x`���2����c#��WG]�J��8
I�Gj&D?�-�<-����>��� �YF1$��7[&�ǐ�Iv)��/�Q�אMgД�
��Y߆`3�-�z�':<���;���r��MӺ��ͨ�]� ��s��*�z�e�Ӧ�������y	�swW�H�|���}�ã7��'��N�����Q�yLe��lTy[�%k�z����r���/j�Gu/h|�s�8�uK�8�^J�C#�,�d
�ݜ��6{½ŧ�����B &�#
?�<��Kz�@���s.�	<�a����42ucz'��;�$���nfި�D�n
�_�b���j����(�ݼ6��{z@�?�+�0������>Q*����D7�䁈L<��Pg��^ ��~Y�1����L�������Q�Z����Rψ�b�&��*����WS�FQj>�)��(V1ն�c�CK��,�?�4]q�:�YPn����5����j��`"0���+�u�ba��V]���M�t�������0էc����1�^Jp���O���]�<@�ߌ�J�6?���a�~zTs�13]�ޖ��f������~�g*�&��ڴOF[Չ�!d^(�@�1_K�ű�8%�,i���Z����mt��v�+L����u�Ѓ:��� ����`�88���B�[����'�Z����?9ί���k3�����&̗�`2���m��+;�]g�K�����=���7"0_�O�z����d�r;��ٞMz�jZ9�O�L�}��+���
BoK�
��k�*���>}����HP�sQ�����ǅ�j�;�H�������t3w�y�sRU�v��#��ze��5�t�o:Qj���qX�"�Ґ�$�%&0J^B8�7|'@�EdK���%�q�g@��/�,�;q��f�/�։����x�MԯS�<��9�j���O���~�3\yt�>հWPv�嚘:��F�aBγn�e��"@,�_�K|��U�h6���pu���t=fK#��ͯ����5;{��8M�v���벾i⠑�)4��R'��=�%M:�\Y��0	aH��Ǟ�i�%݈��%p�P
+8aŦʥƛ�����.Z�a7!�!z��p�Ǒ�G� �8izH���N؎�k�uH��Y؄(�uF����0?C�4�U��o��D��oP��}�hBO�
�LM
�U����g^tJH~�9|�鍘��=G=f�M��J��ydk5�?е'?01�(q*���u��.ɸ�.`�Q��,2N��A���F���뻱d������`*��k`�����Q�-oR�����Og����v��)� �a)��T�h�&�������N��GNL����GA�MJ���eIxaH?\�D8d>B_�EK��p���!S]���>�����W�Lm��l�ɒE��r����˽�Ї�X��!#`