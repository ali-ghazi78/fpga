XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���
����_zі�6�io��2���#�g|d�;����,h��xXC�
`��|��q���PvE�Rk��/L���I�x3|�f�ꉍAJ{�;dY���g���Ú��y�����<�_&�H������ι���?	�_�G �C�( ����[��H�ڡWl% �����s6M\~����R�zU=eE�H(=�5L��a'��2|.s�}����ی�������Qǅ�M�ǒ�LUzZ���O��Y���n��%��9�da,��0�\����a.$a�T������h��S �n( �h5���S��<&��e�׽�`˹��H�{>��O�h��sH��������o��j~��7[�C�8��s��_��q��KJ��I��7�[�� K��꿘����Wv�x���w���o�I���B��������-�?���M��ؒՍʫ5�����+�h$՘�ܱ���rqV�F�"�MT�[�8�WQÃ��nv��^�D�om16ď�Gn����5���_���y��e&��A�b�K��/
bC��p��A���3�;L���z��ھƶ��/��[��)�coC�ݦGњF�6=
�]�K���(+.]��o*��;��鉷y�W��s��,GrϷI'�ڔ��N��h���Z{V`�R��=����/Ym�D���j̍K ��)��$ኣ�����#�W@���W#A:��p��&9ݖ�����'�|s,�`�h>"w�_c���kXlxVHYEB    8096    17801�"�Y ��=��P��}��T�=nM�DhGZ��܉V	�-$X�I'|��}@M$H�@4Za95P+��{��%J9�`#81�!�N���X��ݯ����1E�뢑�:�����S�:��߻=H��p�~=�UH�6��2E�[;��R���ڵ��nn�|�_*V?MC��,�2o*�_�!a���@Q�[C�D�AI��P(�uF�b���We�2Lƈd�����9^Ј۳u�~�&�2��$C�7�Cu��k��PV��%����_V<�B�c��(��7GF�`߲��G�/I��	��C�U#d��j5V���B�{�3
u1���iڑ��䰡���iwP��S�w�<�?�^�R.�K���פ ��:��O���i7�ht����������0���V�����/���۫RJ�o����ߟÝ�a7~��;;SJ��#j�0V[���v"���1tzw�{��T5Fo���
����`v̺�X�k]Cբ�����mM^ ը������`ky�ݼ#�&���=i�qɗ��-σ��8��2̆O�O���� �Q%h�8�O�K]���Vv����=��W��c��/F�H�I���N_���u8�iTوO��!#�I\$�F:�T��?B%"k^��1���c�O�GOf���y҄�}*cj�R�Z��k*���CWe2DS�K#,�T��Ǚ��p ��#r�l{rO@@���R+���%��T� ����9�L�	; $#*@�E�R�T
Nޔu�`UUE�v띵���#c�WJ�/8�v��<gXJw���
�wD��ҋ  ��:��WG�h������V�Q�6_ 7�����暕�]��Gp�gE��W��1>;���:�$JAbg��\�Q�']O��# ^%�,�3�o8N�W�(�a����:��K�y�;C���,F����C8�H쏑�u ��F�\X�LC������׵�An��yF��Ɖ?s8~�}Nr:��w�Ϫ��sg���L �k��J�|�D8��b�R�2��MaG�-Q~�UꞆ�E{�L�ͻ.J���Z�����d����XQB�&G<f����eh�8�__>��Ed�SeJ.��\�N�Nz���'�o��lB������O���9#)�D}���+/g9BD���X�od�!�����(grx�b�K���RBR��E.��MI��u9��5l�vMU�TJ"�G�E����c2rO^��s������1�x�6}�Jl�\{T�f�`v�+Y�c%ԕ���"��9_���������Ưc�a��3F�u��P�e5�����&��F�3t���>�U���alA�~\��ԲZ�v�����H�vCF�tK�s
iQ;-ו]!�Cr/Ur/@@������y�	�K��xC��0����+���Wi�j?����S`��2qƵ�U�Pҏ�$�A&��K�Gd(LT��&�({E_v&!�
:��yz���ڲ���0(�C��	�T�r!�Z�I=�{�v�^�J����ز]Th�� �g����^�z�k�'�6�-����?����E��%4�Fˊ��V_3 JFN����)廬}Ս���n�h��K���,D��!r�N����t5�� ></�����4��B���V#sA���~�r��sqj.�j���
C���.J&�חf��%��☔��˶�����`���Xs�J��P�����$�Y���c��.
^�����NM�۶�gE����V�eU?��(H�]�6/A�����=E���k���)��+���^�X�V�9)Gc��Ե�d#���y�����*՚�x2:�,�f���vN��Tl)Ԝ�d���&�( J5����j�v6E�n��)�1�CP�$$�KY���3��.�4��������K��Mx��;_�d���vߋ?�\�,F�s��PRh��{�]������c�$x~ ��uI$ݺNAH�3O�q8�֣���ZQ-�H��ѷ\�0E
���&����~N�h�k��/��+�(����q �����|��Ng�Xi	��ᄧ4�45�,ޮi��s�!��B`%�Ɂ�'�$[�A�}�&��Z� �_M�VS���� '4My�k^Wà�<\ ���G���Ŀ}H��@��q�	������K�4X�mn�P@:ɹ_����1�/?\4���<�mW�9R�q���`A�yq��Ri7XYE0Wz�!s䔷M�qt�P�Yρ�C�+�^mB��b9E9ߞ2ᨑ��*��3�Yqu�
�P��
�U �|��/�h��</a�Ⱥ�u�O��
ݾ4�Q��tčB�1�B�uWl������h������[�r�ޒ�񹍡hP�=����Ц�1\��$�^�&�(��0�5��G�8�0^��c����܉��w��c߇Jc�O$/����	&�7�����"Z0��F��D
\ۚ@a�q����M�!p:���Ǹa���^����_Q}�s"���� ����4��2_�k�
j��!�ZD�1_?�Y9O��b"2�ֆ`חM����%t*�D0�\@��ȓ��B ;<9�g�Q�Lq��Գ����D��ŝ�UwJr\���s�U
"�v�6�NF�M�o!����(�6��y�!�t��nv�����IdtfA����d�/wғ=�O��_w�3��L�H�GX��C`Fi�����|9�pR>VP�:���
_��]l���K;�W�������ñ�[c�x=c+�	P�[N���G�^׉�V���,_pm�\�����c$�ϯ��z�P��2pz��ۧ�Y��a1���%��r�{�yՆ�8�l���\[]]��x�|lWw�8D)����Q�|Ǳ�z�='�Ԗh�9�����2/�����Q�|�hϋS5��!*,�˲� �}q��Ѵ�=�8V���h���'�CN4[�I�
C^�ɜ�Y�������b4�5K�n'y9��|��8����V½�Y��s��!-��x꒮?
;��af׫��3��4$Lxf[8qy��tO�̓���BҙP�~�|g��&~���a6&��f�����<�$�1@��o�H_G��;����[u���3���'�2{����&�V��y���2�?��߻gQ����f;z��gj�T��Uצ����!��ve�	,�eD�&C(HPS+��Ħb�^�%�p�A`0\�l�_3;��x9�=�+[�/[�zQk���sex!~�� ��g6�'�j-jt�߃��׋�E�=���_Q9D2R���g�%˶���a�J�%͹Զ�A5�8���y��{9���Q�{N>0��Y5g�2��Y�$�&�oY�a�?��}����D�K1~Z3�}�0�2E�.)�HYη��t_�D�π޹�)�h�ٴ���؂��%zG�j;)?U֊\=�o��������_��1{��pa�V"+<��K�����1�Y�ǈ��>�y�4��3�U���Y��
X���U��.rŦ�_wa?�TD�������w��o��l�>m�Qb	T�R[�V��BԢ�U�tG�"o�|1�.�1C�Z��;WYi~%FW�����C7,��,�ϥ��$#����듞O{R����4d3�lP_��-�Ue�PU�1S���y͉�z�؎�fk9�U`k; ���A�����K�*�}�6&��;���������m�׵��+2��E�%@��|���o�[ÚuX�[c�슒��f�)�/틷� 19��i���	�QR�ݳu�Q,�ʁ����$F�M��u:T��d�n���k���F]Y}l������S�^#盉�)ծ�;���*�1�B%s���T�
���vա�_Ԃ�w�3�m��Q<�W�\�?h���0��+�v�[nK9a���lE���%Ϟ-2�28M���0������>$5�4�s�!�0��f0�J���_��5b/���`�h.ɲ��Cn��z�n���j7�5%�.���#�1������*qցva�f�k?�ky^_Y�����Z�Ԉ6�V����"H�̐t��Ys��ul���[,���?�O([=vp�h_{��#~"`���5]�#܈J#�J������Foh�Uo7w)Ȕ����y=�؝Z�lex�PG*F1��b����~�D�$�Y5��k���g��TX�CԲ�g	K����	��������:����!����&X�6�a�ێ�yި�*鑾N�^ߘB%��|�܆`�+���Y[n�K�t�=C�E:�����o�dx��u58�6Y5�4gD�@��Y��b��k���w�նG�j>��˄��kϢ:|�F�,���N,�5��T��oxY�cD|�X,]\�� �c��iIol=(��A����Q��h���Ʋ{�186���Y��iɔ�O*�6]VV���������U������i���X�X�/���৤�l��W,Ml��;l�c����7Î-�>�{t�;�K�����9Sp��}��-����'{��q!�/2O��\��!B~�dM��D��� h��$`��B:��="ڟm��� s��!^�O`�T�cҭ�%`�){������[��uH����NZ{iL�@��]�K���.�_(���{i��(T�ǁ(����Q�5Y+����Z�ԉ�xr)tZ�������y3Ns�NV�����Ci��u"k��eFc�oG\6�??z�RG�0z�/LNnE��z�,�(�U]�ݱ@��ف_���
�%8���SUM�wr �1�&�o�84A��~��~&�P`D���m�#ᆬs�S�<8�x��7��=CG]�k����E�4�sKU-G
=C'�6��1��B72i�����TVB~b�i�0�N����զ��Y��� +�<L5M����(�C�c�WH�e��;�)�v��ݟ{BF&��r-�m; 1��������#z�KKI�*+�/������"�(>ukZ)P6'I�@�<˃QJO��&�<C	bн��\T���^��[A�pL楼t<�|�j��d��x����'���V���h�*�EQ��=��D�M�k\/���� %�C[-G�yT�5⏏�D �5�_�lis�<���:F���,�iR����8n�D[$ɔ�
Hi4���tP��y튭9)���d��3�J���6*LC<k������S�%"ǧW�~Ѿ�ě�O�b�,�|��r��A��_>Ԃ�-�[���C�?�Vg�7Q�?<!��a�$�&������i~1ߦ�\������K`�2�b�K_q�c��������İ�@��� �=!�x[^��+���7G�y���9��4BJ�a��-|�G��ɞx¬|N&��1~��,̲��3�`��J��Ǐ�l%rQ��⸕6\���y6�H���+��������).4n���AoE۷"��)�IC��!�� E��'R;CX�~���?j�6yd(tǣܩ�w?�Z祰Op$�D+���T]�k2q�����.i��rP���O�8\)�+���'�M`���A�s��
��h�#9����J$����aR�˓�$����͖2ǒ+8ϲ�����nAI*@�_Я��<VnĚ��h�\��m��\B,�g�+�fY��+x�`E�<ͼ��H�!a� "���ݶ�#N�nT��7�{�n�L�à&�:g���ī��,���b	�4����~�!r�;f��]*h'4�"_�r
X 2@ZF
0r��p>#�5��I�H$hۂ��WG��e�P�)2H!���:���\��m��' ��}<�b]cx#��xWE��6G"~�q�r�Z���-��:,� wb�W��TrC��
~����ʌ�A7���D�D�G�0�%��e�w7��<����-�#�s7��G��kD�X.�P.KVW~�m:Br	D�W��rw͂��m��z�ڍ�s�C`��O������q*��]�M��1�L̴��t7M��u�O���ɵ("N���