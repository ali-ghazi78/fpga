XlxV65EB    a04b    1c60u���R1�̇�?�C8�^�W��/Ba�V�7���%����7�w�^��h�f���iW������I������yz%����=���;��*r��8���+�{��]�bg�]�3�PE6F�8R�V��C,��U���M�+L��)O���o�g/)->��j&��3c�?��4WA��V\��� �N��w+�z��ՉC���I������� X�p����p�m�Ο�Q#߳Z�]t@S^�噐C�`_G=������A�\�e�x-fc��<A���KbѤ���y�7�<��B�����Е�O�%e8S������1L�~�|�v�k�',
x��$�C&�j�1�5�Ze.9���P��v���Z��h���Ӌ�%:����#^@�� �P�"¿/i0�����`��ƫ�*ײa�H�>fUa�F%z����b>�(@Z�`��1��+�*N��o�ϒ�~VaVk��JzQ��ƭ�������-��!�X�!t:���=�����Z9�>�d15�۲2i����f*Nz���c {QZ�2�W�v�#<�("8��_��z�(1_JdK|5�^x��
��x��D.W
�C>�A �j��7k�oF	u���ЖG�#)��G�a�z�,k�S@�:�ꣵ�va<�o���˥&��u�Z~��:8Pe�x7�% !)�\<~�m��5�D�I��=�m򎊑 �t�Bc�UWu0�,Q����\$�N�F��Amz� �󯵒�3��5���Dv73��gc��v�V#%�D<1/v�w2�/�<��!jͭ�+ɐ�V��>���C��cR&�&%Ԭ�V^�I���%��������|)��Na�=Fy�.�24f��;�8N}~��dbY�o��%?�.u�oY����1��j[j��	����ذ'�L�!zAp�yԁ�6�Gт���~�ޕ)�a�\}� z��K�ʝZ��K����H���o���+��LM�zO�iPY�9{Or���b#����b
@1,��9�A������`�/�(�;)�ݳ?~	�L^j�-h?��.���Jy�������4U�	@~�6�ge'[I�sz�Jl��:��q~T:�ڎ�40�!GL�t��2��$���~2[8����M������i������bM���p�%��Z��u����	�f�)ME��$4��qYn��9aݬ��}>��{툡�P}�!~� �#T��(���=:}�'�����I:G��B����a�>���G͔]����s��5���c����=o���� ���E�6#V�Wt�Ā#%�,]ώ2�����i>�s��k�������Mc@�_��/C�6��5b�U��^���r���㪶V��Z�wSZ[S�$�QK��ľ�b���g�@�7&TB���m���e94Dh��o'|0�ceP������U���2;=��X3�/��^hf�m�ג����jY/�}��� m]h��rl)Mv��\����g�	����S��)���j���Y�h�,�}M�:��Ћ0�8~a�fB��8�F;;��Wo|D��m%�f6I��9��*��������(�a�E��}�ۍ��T~9f�ś._�>3���H �|��M/m���+ Ȫ��Tt�Z��O��/�&���kf���"��7�޾XR��<��z�l��/�"�`�P��ҔW7*#J���p����H�b�ߏ�5_*^�'%x�X�C��EcE�������z��Uڄ �(o'��IdX��ڗ�p)@���TD��U!�Jo:���+�]jH}J�R�������R7Cn�O��s� ���Vb�U�)Yb�W�����
��%J�Ѝ]���=G����g-�S)�"���`�����m8�{R�0�x2��
;#���l�ᖭس򶡳ԵR,�;�5d�a�&��g0����G��.���^�dnz�M;<���Z�3��$��0]C�^����p}ց����&��m�.�z0�d��k�!�I+\W,
3
��=ΜGԶ���#TV��a�RT�@�E �ؾ��2���=m,������Z9>���_�ʙ�Rr�a�*��49����ߛ{`��^7-� r�,H���r�P��(��'x��ʔ!�؆��q�
UDLs`�&���M���>}'��T�D���d����D��)�W�w�+t�Չ4�B��)��+k�/FZ�t�~z�}��p>e�*sT����G����"w�`�����eS����Q�Wi�A f��)?+Z�U��%�4|qX���!�]�C��1�F���O�b�����{��\��(�g5Y h�{8w][2a׈T�w��\CO۳�ɂ�H�l-���긯����'2<�fE��
���=	�J�~�� %�g�� ���cI x��|���#�g�P�*��@�nƊ|�m7��R��p�@dr��R�TQE�̍ǋSC����6���J��/��!�V�F [z��k���K�3�	!�Ւ;o���Nî�� ,𒠹5Ə��4Mc!,�Wk(��i�7��񶽄p��Ӄ(Xl�}��Y��m��� �ݼ�S!���e����ȷ�X�	�S�2�t�Y:��P�;нA͛�9��	ӭ���W:��KW(�lW��� "O �f.k=��P�Ĺ*�G�1�g
��y+)��������!�����}ߡ�B���T�'x��p/��l�8��]g����>�+�e.N�(>���RJ�A����v �R��WO�^Ԁ��.��9*\#"؝!ӶQP{gP"ƋL�O��2��ii���=�6sy6��/�4�+��q�OSV���G(���OA:Q�P�:Z�Y2`�b��q߆K���7�=Y��z��䷵8y�rx=ˠp�2� 3�f���I���	�9�(�8P���_���v_
v�x5����FA��ҫr��-��_��<���ȍ�c �v��1��x=K�4�oy��U��Eˏ��Jy�b��n�uSc������-8�#�R��N�f��ޖ��x�f�~�o=7υ�w�j�;�����G�p0����#,&�J����ςR&a���Ȫ���ե�f�ΤT��*^j��]C�@g���]��O�U0�I`jm�F*0݆�NnC�"Jms6]��|��[��ib�v�~�v�P�9!Q�v�\�QW��8�丙�� )5��Ag)gH1�kK}ʷOb��Qd��ܒ�ȸ�1AS�m��zL[��q��ʞb��vL�`^A��+ �єlV�*Y?z�N3�m���Ǩi͡�����y�U�;��@jܔ���-�����/UW�+)�'�}�7&C�����>P��s�4.�!S��ޣ�q�sn[��p������:T?jF���������$ŉ����㳺�Ÿ � �Ġlޅ��F�}X�l�����W���Q�� 
���N^���֯h�O��B��<�X#ҐC���F����F��qk'D�P��%Y�:&�D�]�t�q�an�y�P��Q:!����/ w�!J��sK������+���7j�4��~P!��m�#sL���5��U��qc��Ι�й6U�Бes Mc�{&_x��mC�D�&�萙]³�"ɊKS�NR{���������C�����u��c���%��(��ʓ@�7Yt��"̥v��Toˠ���L��6v�e��P���~��z��!x�Siq�n�?g��
�J�y ��e*�h �W"���pMz���f���	�������g�l{)���m5G�|DfJ�x���(�9H��TT-Sr��5��O�V?D��Fb �Z��5Z�  O)g	Wp�~h����C��s/v䧽���i3�S�V���~�"�2�v�xs�b�����cR�ت/VF�Ig�-���NdV�\]��:�^��|  �х����j��i�c�X�y���Y��J�\v�\}}���T������(Z�x�^	�����l|�`�΢п[� t���Y��,������n�Q���#��H����A`-(a�X������	�t��<� \�Eřg+���|�~��'�%���7*Kؽ�?Y�-Ofu�l7�Չ���� d�qo���׵��-������dbW�Dw���2�xA���5Y�X��mBU�W�k�������q�m����Ǘ{h|u�t���	b����N���g{7���:̯/�$�O�]�7�Jӕ%-F,�-K+�3$I��,�>c����ua��|}cE�9����o�N_��û�CGŧ�3̑�D���^L�(�����I_����	yA�Y/�J�6'�z�������(�ZU�=�G.�+��$��Y;���I�rр�!�1C����r����O��'C�u�MYzvr�lr_�y��f �,�ae�F�S�z�?�p=�Ȥ//�P�3���Q#�����Ý�E_��l��,�|�=���H!�ۇ�ò�4�L��S>����-ƪ�<nN�HBM��S��eG�S��	v^��`��ά9h�h�==f��z|E�v�<���5QO��rM��HB��G�M�n�*�O��.rR{�� VTvƊEt4�8&G$�so�_#�kZ!���?� �X�!L�"��B�?^S�fN�)�,3�����	��������l�H����GJ����b�V���֏��¢��!��o���U�7�Sb��{Gy&��l�j�޷{b@K1}���E壕4=f���3��<Rf��(�;������=J�	1X� ��������d^�,�	�,T�:�V@/s�۪�AR(SEu��CJw���d��h+�=�2TY�U�������bA�ߌ����ZfN�.V�,���f�_ڧP�,<���;w�N��Os��uS�<�ƻ��;s�<���Q�V�n����,\��-yn��Q�;)��_y�{H|��9Ŷ�8�&\��#�-X�rJ���{T�i�i@͆*b�R=�aM���:�$��r�VSk(���<n|#ޕ���GA���� {�uO�412��΍��(��
D3��I������>�|bܴҁ�B���و ]Iǘx��A�zUĘ!1�n����j����������ai�<"W+Nz�+@���/�MB
�Ӌ������#r\�)�k�C]O�y�HIŊ��ig��Jt��*����G/��q�<%�tÙ���*� +�zKD�V_����N�@x��@��`�+`�l��fO��9�έ�px�}�؛��s�СɫUl��/VdӗM`����%ѪN�%���za��8�#���(�![/��v�Va��7��,"c���*�����5|�S�"���l�(�!�(�{p�9�კ%�z=R wG��)a��ɟI���Z��L����?x�����
�̼�/�u�i��I���wq~��V�5�����|�[��I�)�S����Q���2R�E&����[]t$�z��c���3[�8���o��y��u��E^K���JGs�<�ML#�XGO��V��H֭K���l�D^��o�;�˿qL"���o��v�l��L�~�r]ƘB��+����T�ڣC��82h�:�dN�	��̟\ǅ.UeH��,�.>�-`Z���l��ބ�X'^N`��*�#H�5�c�ٖ�N!�]&�{����A�[�vd�ULE��1X���OAR�9!!��)ީW�~��)#�â<���愹]N鉉��<��z��Ct_�S8�&<Nv����G��x�:-^z��Q��J�P!0j �kT{
�7�MN����7}���܎֯)U�`~��ٓ�bQ>Ϣ8��i�� �F	��t�4
��sv���x���\��eǑDh����;b_@�\����������L����pL<����_ ��x���C�vӹ����#��6�/D�X|�v�(C�����!�[+
�����f� �w�rn���7���T��1;����^��b���`*�DM��'b㑨: �c6�� ��V�4tI6�e]k�2�y�~�ՙ��)B��L�}j����h�&����?%S�.��������3UĨ|���YxQyC*F�+�K5�����Wv)�g
A���t�1K���;�����~�t{Ft]
���iz𠚂j��e܀>�_ԋ�&�������>�I6��M�s`�,t��*G��Ш���MX������ʔ��OU$�"�'n'\� � :X���������8��,#�?�O�b�?����ھ�%�,�0�t��= h�D����7�?"�ꢻ��4Y�nVL���"�G�.U�`�jS��=jp$�磾��9����l�ze��]mL��"�ݯ����'�h|�O��1ddh����5L��.2��Qw��rj.LB�/�x[��X��	+��{F���7w���[hˆUB���`]a��h6���)�	����5�T�gpm@�%"�\���f�VպIKG��[��-_sB*f��+���/�*ט7i���
�����a�ӥ��˖[»t� ︁�y� ���B�P]����M�S���{SrЀ��I�@3\��Z���c|��r�y���a�G_|�\�&,]pR&k���¿���=�f���`/�6�@�#j���hG�2 �!6��L_������Z�!�yv`�}�ބ��[�H�y
�FZ������jM��hg������P�>=�N;�7?^c�[m~�JN��U�K��+W�Xֳ��{�e��!��p�jb��탆����ϛ�!�K�p_�3��!jǁ		F���^_׷
F���[P�9#���������L2Hm
��w#m^~�����Xe�VF�'+�R�QR�T{Z���pм~ߪ)ka��p�R������Z����`�i���t�Da!�SP)�.`fAg�xz=�lC+nv`V�'m���N���/���B@��H5I�f�A��1��������rR�Gi��M7�n@�5�V!6BTz��v�+�;�*:,�����C	~KQ�>Hk%sRdg�� ��Z�Ą;�N:�Ϧܼ+J��YH�O�pN.�7�J���ȫ�oI�m��|�y��r:��@�&e�"E( ����HP�!����P#�����6���EH^�L�3 @���5��a�z;g����p9���v(v����j>l�bDd�c�����og�H3�F�q�q+%f>;�@