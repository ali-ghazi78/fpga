XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���q�b�)g�ty���HW��s-�:��C�aI��('N�����ac�x ] �^C�/����cf��ܤ`D�dJU����:�^��|�d
W�.*a�����<p������{���m��'	���@���'3��,s�=z�q�3pC4��t�[�Zq�����q���	R�qs;�q+&O�$[ǿS֙ ��ioK�h�S@4Q�Qt�ԇ[��t���mvQp-0�곆xlG���ڪ$����3F���
J=oSv���)�� �J ��qI�Nj�^no\�vZ�3�����|��g"���im��a��΂7�;��'����>�D���	���2r0�����,X\%����{u��3�UK�V\:�_w�N�~�e���J��&�E�2��s�h��Z���p��\�-���to��Z{�|�6ռ1��!�f���j�)�)����O���'�E�J�a��\���RfJ�hQ���Sg�2�*!"���j�y��s��\��$.��;9 ��|����q�5������g����[�O�S�4�:�ÁF�E��)Ĵ��f��BPOA�B���Np�1
���}Ym�cS�b�G2���ö>b����������d��<`�_�q,���X_��~�ܖ�$t��ʚ��q`�6;'����[��Nd�P�);�u�_�s�
Pڌ(jhX� ��\,pb�p��<�uNS|`�NvNF�'P\�p�Q1�'�;��Uq|�Ԛ ��=���4��+���e?>:�3U�;�ͥ�XlxVHYEB    50a0    13b0����d(�J����p�֋����c=��m���.v}n]��� ���u!ۖ� 0���}8��S��sY6�����cu�`0e*5(9��(|J�b��Zf@�J"(�Ѐ~�j�6@���<�Or4�)��OJ��Y� F+AYfR��\��Y�A��"|����+�z2�ZzHhEjc�P���˒~�o�ۚ��'|�xL+�5�("��֊��ѱSg�	|����泤:�	 �F����U5�-@�A[�Vʩ��}�LYL��BHG\B.9%��Қ��'�/:�B��A�4+����k`$�%�B��<}��j0[��]}3�e/���NhU�6a2�X����D���o+E��e���qv�U ���>W�Wc�8�{o��M	���Nxۈ��]'��,D��RQ��m-Z��7VZ���"'��4jOm����"J�%ҏ�q���r3�?��އ1G�lD�3�J�� ��e+M.����C�7|_T�C-B{5��;������z�f�81,���:�5��9r�����F���7������d��l�ۧ.5�u'��v4c��X��ͪ'���/��8sf�;l�Ls�����j����ā��d����o��3 N���*��������4+�kT��9�2�TO#��\��F�V��~�����덎3�h�Ϟ���$�H%fftQ]O��Bq�!̝�Z����P�~�^k-�P�$N���:��ǎ��U���«c-;t
��V�b��LG�|�q���
��91j5�� +,�_�cj��<;��r��g�����q�&�Ъ�'O���q�� w֙�>�mw� �U.�Y����^�E7_�SY�Q��1�г�
@G��[��T�D�/�@�'�R�+A�B"(��φ$UT��͗��/q��z�r�<���4!�_s2f ���M��YW�u�Ûŷ��i����L.���Gd�R0��=9G)S#3'�Vr�%]oER�����JJu�S�[&�@"`�B�A�s� �����TK�C�@��� Q���Q4�@3�[1��xC9���c�r��5��+���S�3��c�P�Sg9�l�]�U��"cܛ�͐�i�ػ��j�2�[�^�����ﵵ������g;���oP5��ޓ�ΞX�]�t�(vC7��G�ۼ`���eA6��F���n�K5vl!����(8�q%�x2��_9f2�C�ye���K��ԵA��J���D��R��d����Y������u>Ct��N�I@�]�g=�Z��N#X�Ղ��V��"��f@(�6*�L�F�Ц]l&�v9�ɒ,&~�n��.�|x�� ��]���䀩<&�Fķ�Ir�/K��,�naf(���Ia��GF�ŪS�틺?sm尳���\ɿp�|m!��V��Y^�a2Yx ҷ�yI0�.�EhX�z��~�J��{�Y=n�D��Ql�wPm>4ˆ�T*��GC�=��Z��w�Y��+�{��._���h�d��e��@yMZ�#��G)�]���$R�3}H��қ%T�2�u�R��Bv���i��]�>0p)R3�⑆�5Z������a;w���#�u�^W~�i|�dOI�I�GA����5���q�H�we����#*N�]���m�v;�Nnӝ�{Ȣ?�'g�������	�}@XW佰�!��[o$)��|;��u������A!A���NKn��Կ�F d���mK8��>)L{��%Zs2���G@fys�zj�����7�-�g:��`B�e��(pR��l��H{��� � K���UI}�*�7����n.��<��0x����O���'I=\C��$be3#�f�osL��]��a�䧷����-8�����zjpƄNv,�ֱ��?>����hb��h�AW��)Y�nk�b�A��~<Y�����YjM�8
@,�,+PӨ��=α9�ZC��`�lwSs�ϑ��Mh]\�S��x�l�/h�C @��=L	A��	ŏAP[�)֥��G�OKd?ٛ5�aK�ڏ1�b������'�؞@��Q��n#�˂e��82�;<c�Q��@Pm)J�B�r꫊��6�������z�sf����kux\�2[��|yR���g�3���W���?�|�#���>�&ف�?�\c�b�#�������Y�㽞��^&��<N����Ũ�����MPH�	�:��ڑ�$��\yh�����ǆǁ�I"����8�B���dE��!� S�L���ʸ$����s�W1�>��m�����{���1D�C7����:�BE�tCYS�	.���`�f��<�G��P⠼�^�kD�Y}5R�o�kae��GvJ�����Jea���i����.�Y0Zh�zV`���RĶB�C'��}_�ݼ~�_����[��^F�#hUD����;�s�	��M���?��ff��P	���
v�e�-Fx ��c����/��7�~��א�~c��<����v�==ae���&�(�7���94��Ų2Ң�����c��g�7v�b�!#�@u��D`Mr���ݏ���8$�g?��!qij=>M=<Ɯ�wLwɻ7l'��V�L
I���v����Z��A<;��:��iqy�X������2���]�7�;�#}�=���$��K�N�Yi���.�8I��e��RK|�6���펈�o�����
a�i��������~l��g�s��qGU�+�>���S ����k����ZT�PW]���f	���q"�qbJٶ��k��w�w^��5re��?����zg��m1� .L��m8����L�w!��Ń^�a�?w.�m����.�M�@���z[sX�V]�>_`�
Ij�Z@���!xvHX+i����ZK�
�Q�[�6�Na޳���X�7��U"b�qv��6�W���I@-Ry^�B�<���^Hu���x)S0������'����Q�c����Q_��B���n}i�z<��,ݘ��w����5�xR��U���,c�̛��/��{ >�������Hol^$^G�jh��� P;����1H̡�.�P������U���7�C&�� �ؔ��w@p)�-ӑ /��R��<ӣ��G�ta�.a�x%NRY�ո2Hj�p�`�W�&��_>%R��sT����)�b�L�~��(zW*A����Iq��M;ؙ&�H���^A":Ѿ��l���2�*r|�'���L��^�Z+��3��0�cF����D�� {�,��^d��;�'PE]hÿ�x�=
�5��%��`�H��������~�FE��G�(C�9*�����C��9U�a�,/j�����
�6�&/=�B���Q��qT��
��n��8|4�%�4��XH��ZW��Q�H�ԓ
V �����r�T���>@Ŧ�UN�ۧ'������s_��D��,�~$�k���k��{���eLs�T����d�'HT�����`���g��[�̰�'[�!�3�m�P;�t4㛦K_@}������ &�����3 e��`��ӎV�	�;s�����̨X�C�L��K�b�hj�v�Mk>���'n�P�,�4��٥�)���3�kB��E
�����h+h�L~E;w~�EKG��6�ˢ�0��yK�����(�h���Q"�+�H�N`���8�9Qu����1MXy3��>�x�M��9r �x\��N���#�qĄ縁0�j�m����/��}�q(�V�fVX�f y]|T�� 1+����,�0x/����`� ?�B� �ô��X���m��r/e�%T~>V�5�^��/�1|,���k�vg�[�YԀi!�G�5l�E��ж���,���)F�`�0 �5'K!��Y��kyX$�+c^g�z��iÒ����6D�J�A�KPn�_���9��)ܦ8p��$T�"�2��S��|O�dn�10z�:j�M�р��o�9z����![�� �Y
:Q��@��C��	^�Lc9U���V,8�^�9e��[g�Rh`��t��B1�TW�F���-}O�j�O��������yc�H�@J�Ʊ�:�YB*�/���,�\[�����F���<���puBu�ʦ, Z!�,m�T��Z���Jz�fޥ��x��C��vjȡ_ub��!�5�`���x��sД��L����������V�n���A �ۓ{⮦"��)����fk�Z(�����XQ�Cs��]�ΆՐ賛���Ѳ,+���L|�w�)3?$�#��閟P�CB��@4�ė7���h���mR-N�g]��|�!��=�<v��^�!϶F�>,m��M^-b�kF�����	�����)<(0�ڃm�_�h/X�lj��Q&��@�������:�B-�\��?�[��W�[�R}�B����0��R�C�T�{����F����W,�͐���.��>L��g��	�3�]�~E��i�����d�Qd^��a?��T�m�g�B���-R3 �t����d(P������-���w���2�Ev��h���5Ѳ��b#�Q'�c7�ȴE�F�t�Ѓ>#g�ۧ�k-�����YΊ��߻5����dr��9����|��7�E5��q�dյ�lԹ��_�⿋�[�j�LҰ�1��sGV��Y,Dg�<����c�6�n|ggf�� 8�����;��*p�S]��eRl�u����$ь��[u)��v�OX�I�-u�3T/.��P����]�]p��H�չR!����08qVU�\�0,m����S�f��X)dՓc�BHD��^�M�I̿�\��U�����@�Q$)��)SM�{�N)���r++P2������?��� ���Xy�1��KM�A52���~�l�ǆ�<y�����q���+[������;9V� �.�%it�7xT��DOON