XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���a��O����f�ԲC�b�:{m�h¯iR	�7�n��^�>OF�O��0I)����Q2X	�Xm�t�q�S�Y@��PVl([�(���
����\�ؗ�i�+C�`I7���@bc�#��a����#��7�`��L./Cton��/�W�A�	i$}�n���jq���� -�d���Tl�����JbkXX�q
�ǫh��sh�-	Y��6S��+(�yF��T����@j
�#!B�k,���R3oC&ȃ�)�M�[�*O�59��� i�:j}ߡtff/}Ϋ��{3�pbz����i��K�U�G)�8��Vj�[�d�B��%���&����4�3��VƆ86�ʒ(��9�ߢ�-�˝���Ǭ,��X�L��F����+T7:.M:���̨G�zO;��с��V��;�L��J�q�~�[Z�o*ְ:�p�)T�Y�ʊ>����n"����`
��/�-2�+tA*	�K̨V��H3�!���!�	�n�>5w�0�e�'�(��W@{*�L*޵�\�8�| �Ẏq8�L?�S�D�_Ξ��+����\��+�Hdҁ\c+W��!@�G8�,D�ؔ�N���؇Q'k�r9Q���9��m��Ȑ��a]rT�k��2
/�xAß��	�����P^we�Q�\=���lr�\�u�ӯ�jxY�c{BF�������\�k���9���ؚ2����V�F.7�H����eiԬk��#m�y��g�đr��"AV�j�f<ė/�o���XlxVHYEB    6a5f    1320�ڎ�7k�r�HH9͔K��.䮒��˭���G.|Js�ῇ��h�G���+�m���&�;�]iE�!�9��Z��:�e'^Q^����t��`[�6%��8VJ#`�Z�i�!�-�H��Hpɟ8��a9NS`w��-N�V�R��Թzo���N�]!ڀ�>�6p��U��d
�^zC~O�j�j��f:�X�4\�h�Hɧ�O�E0�]���E��`�o��K��nC��S��Z��e�����=��_捚�nިL�}��+��T���b���"�G�k)§����BrTcD���Ľ���پ��>og��ه~$�\��b���u���M�ՒY����P�+�Lf��D"(��#�6�s
�!zQ�nz���Ah+���8�g�i�d��%{83Q�#y1�Tݠ�X

�5�3�eJ��<��m��Ή���jĒ��;�g���:r��0>Y�n��t�~�|@���}f�h2G���b.��@��E�����^rD�����y(�p<�� �!G�ٻ�E��$>����0�"K��ʦ��}�cu*�^�ަ�n��N�]m�����8C��ߍSF�+f�]�A�־z5��	dSbB��r����]�I���Q�FP�b�v�:� B��y �:�'~��=>jtK�E�R��#蹒��N���'z��K�%3W  ���tc��(!�����(�i7�-/'_�;	�x�H�a5�A�hv�H�pZ�lPX�)��y=b�W�zq��KZ�-��~0�y��,��pA�-������Z ���ݘ1_�ˍ8����L���������>l<��J� J�"��D�:K�i�Ϩ��aQ�U����U�х���P�3Q�G�g���~��m�7���#����7��� Q�f�9^4y�4��ep4�ަ'륝k#4�#����ae��sD��`y)9b��Q*�r�'i 2?�������C��^[�2�B}%\e�~�>��yBS�a�?%7+>\e�8Q�>!T_W�7u$=' `(`|�ʆ�c�p���L3�kH�0��^�d?Ѹ�|e��d՜�Qf��8���U��Y;��i����`��'�\�z�xaz[B@,s�!�pT�>G-tE`��B!�BP��a4��F��Ty�;a��5r�D�L}#v�c5`��khf`������� 3և78Mq�' _lpݫ�d}ٔ �Y�#yG��.h��?��U=wn��&�98p��$���h��O�Aq0�҄��]�LI ��(�M
��;�����%�x��)��|5?s�����A<��4�;l���\�N���q^�NLjj�;3�WRX���f��d�lk�r������2��.I�
^�#G��U����-�8o�܍'��r�:F�Q;�$v��ݨV����G��I=��,2)���pP�A���Mp�L'N#���p�"��݈�ۆ�=@
.~�n��F+��?���v8��"9��@ ���yL7??B�o�u�lEb��{�����}�K�����W.Ӥ>eVQU���N~E��n�f���T>א1����K������^/{ ]�!FYx���Y��R��*���EG`;��� �������,,��u��d5�}��H;�,�vh��ߵ��2�F��`��W��k���8.(b
�̮=�� G6�yx:7����+�\�P�m�<Uʖ�h�7��=RBy���Ά�PO{ �c5l%��D������J���P-����#а�g¶��X�i��8�i��=��/11l�~C���`���i�~�>��1ci�� M��]t��NIu�G�%nޞ{�s�o3)�|i�QE� w��GSB8�����')2�m0�5�0�ܼDIXl�B9�7h89�	����`(�U�D��jV��+,��5�4�q;x�+۳�R���_~n��N�	ư�0XsQf�>�ה�U���#^$��9�Y��W7m�DzFly��r�p�k龎[Д Q��*�Q_,A��O0���P(g��"K={<ڭ��֤۠S/ܽb)�����#�������T���,�Pa�ь*���D]J	���.xl��{q��g��'O�7r����	ϛ�}`�*��B5F8��BÉI����Ղ�`�X�]��޳���e/�qf�Z$X`�$k�lj{�i�Zl��zDp�6��~�=��J�>�жh��÷�_��%��Dř��Y�ם����c���%��p���&�Ȗ���v��j0��e�K�b8XbU��%	a$�GY{.���k8��mqk�C0��C+��t��$�T�FT]9��g������\����
�kn'������13������D_��%\G�G*�n+%Ϝ�*~�z𹇠I��Fj��:Ho0�ɄԻ�1q��͑o�_�������+`ga�f}6F1��(� ���8�^l���3I���n ��1ę���Cw/ι1�88�]��N�!�����+�(X.��g�I�4:8������>�"8�.��a�k�-D�/��2��m�;��/)��_�}��Z���a�0��B@`.����w7W��^Lmj3_A(�<#��`%Y���t��de���?|�(e�D�^"�>M-؋fR[�R`��%gw�����DdAD�o4�YE��m�,�\�ɖ�@e���'N:�;|�ߘ1S�v�xaR�~U���Dn��N1�^�(C��jC�f��`#W�K���ѷ[��A����<�]�w`�/A��R����d%���>�eX3$�v��g����*�0� f�rɪډUhZ�Z���VD|)���D!�d0���vP/� {	K��HG� �-�>��o.Yp}�!*��/�$���`=2��]Aҝ�lB�'����:fM��.��
��9��{�;��@����OQ^��1�*��V�Q��Z���%v���
� ��!�����ڂ&��9|7��?)�_o�(w�=�;�����)}�R|N��iC�W]��@W+:�ٓ���E{����1�(TJY#��| �����f�ٮ�}s��;�!�	�qX��\�3a�k�Zo�� �ӽ	�)��^2���0fFI��h� :��o`�$<��6��Ao�t����lF_LO�XT4���c�B��\'�v�zf�������
�a�}���\��5��O��>+O7|�V��Ŭi�W����$F7A���q�⟉��%�?]o��N��Q�Ɨ��.����g	�7�Ā�	S��`+�X��;�8Vr� H��T�W{������������Y��=�iY�����rS�l�̉�g�� ��*�Bn1���][�WH�˖O�v����Z5I�4��cs�)�T��d.���mV�}ŨH���[�qX�psyU���k�1�+�D.��ƭ��B6�c�a)�$�c��I�8��������:Do�z0�R�.�b�l4�{�.0��i@�v!�{�K�-i���z{�v9OV9�qa�Z�:S:@���ݜ(�� ���ba��:��㜙���b��Kn�D��O��8�� �@��/��ۿ�ɻ��	�^���z�tM�;<ER.�ന��JP\��3�%+���Xzh��1�--[]�Q�u�fX,�1!��m�sd�zN%��oI^�NͣZ�����Vhz]��zz>Z�4(2U(��Ʉ�����sS{ϑ�rV�#�~��?B�\�6��6�mB\��@��<j��z��6$Tu)_z{�`�P|��Ԏ���v�h���~�@��E?I��(���2MO�pAH2��"錆YIR_��F�Rf�
���������w�O*�uJ��n��0J�t�:XQ�.�����R@h�w)hg�x���~�m�͂�A�%�R�Иi�+�R��i������{��m�-3���|��j�����v�~�R�
#�؃2jJ��7��ʅ��5��7�Sd�	 }`�
O0ί�H:���beƄ?��CYz�>{��)����gP��!c���e/TU�Vr���u5�6U.l�g�mN5�]܏�E����G��M�@ĕ��Ï1��C�7�F�,F���5��"w!���~q����������F�L`G3�e@�4Q�b�2/�	���n�%6��<�K}3ۦ�#��G="�ִ
\Yue�2��Ѭ�*f����J�FG{�=��j!��� ��$f;'0����wh��Õ^�Ɉ����I�(=�U""�|��77zs��Mʮ�n���ܢV����{72 ����vW�>4��S��t{�յu��hs
&+�t�A���,�=g�M�I���UZ���(�q�
�5��県�#j Y^��ۙb���g��XlA��G��r�������i)@���	�F�r���)�u���D?�����]s10UR��5�G����*����w�^~0����!�g!{HG��IO(�1Ϸ8�'=~�� 76�K���$&�a��C��'���HT�Ѧ'gSC�d3���\(h,��Bm]���kq�K�cQC���<���Є�5�9�����m!��~Iq��G�-ԑN6J60��� c�N�Y9��iX��a��G;��]�Er��2 �	����\e(�k��3aƊ�j��wH,����R�j_�x��9��0 }�_i*��=����9����]��N~��t�����j/_3��]��6B�[G��l[�NB��4t"����@ݳ���Pp1n� +Z���hOQ�R41�N�4| ��SAUJ����;f�����#�^��Y�J���8#3�����4=�F���K.�#�\�aqfڽ.�MO�Na�Q�P���4nm�ʲy��e�A� ��^Ko�09!x:ǿ�GIu