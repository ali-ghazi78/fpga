XlxV65EB    509f    13b0.��R��tB�@i3C�a؈����hW#[6�^o�5������Ćm<AW�J����'���B؆|OLC����^q�֕�7M�[`�����e����"�b���"��^��G���\��qC�@wK;Ҙ��r>��"�e�q16蟭$����ՂD�`}����
ףp�j\�_s�5u���}���
�|5H0�@b^��VEh��
�/�.E&�m����Uu���A�?`O� ��;�ˤ�{i��-2;bG��1�g���r��8x��M��<�z���~���'J��*.�bLO�kkt)d��R�K%{7w�B�4�˯�U4FppB�N����J'h9���U������c������Rj�f�>ۅ
x$�������B����!F(h1�*=haPTc?��A�m��1��W����i?jrh��<�3ߦ��qҥ����1��"��0#:ncB��Βc����Ku����2�+~�O�_ջNʗq	�W뱏�b����J����-�#�@�Ͳ-���<�c�y7��hG�<ٷ�y8�^�~,�󈘦�ʠ6g醊�*dث�&E�Q�"��s��3��7��i����i�0�K�:C8�uq�d�F;�9��L��2�,��*<a�{qՊ5��q��VDY��hɕ'�f�� :���ג,����M��d�@\F�CaY�^�M����6b��&ⵀc���5ݻ�i���c+"af-��?��s�gh��6z�3"�S;c��DylY��OG��H���M���ŦV)`U}v��2Q�h�5�%�7�Ф:�z(�2$����Q_G	追c�A�oV�g��ps�c���wA1�x�x�H�!��Ssq^�#�:����Q�(�?����R�Y����I�-����z獵_E�F��U�y������`��]�ne}Q}����H��G-�,�ȜF�U�ކS��^#0��d�T���$�� <�Q��Sf��u�+��&�:�R��#亟�`2�d]���u�����.I�=�z*����L�Y'�=B~]�T��}n.urρ��,��<� ۺ���Q�������4�*�:S�)hQ*�w�@.�ث����E����Ř��'����'�r��#�F��c8$EwM�i�G1	��Μ��b���0���*ՒU�-e�>�Ff��8q�Xn+�����;��r㈰L�<�O!��H�������%�{|�Puʿma#�1J���HB]i��M�V�cfn���Ir��ї���jG	�C1�g�����ɔ�}�94�	�BF\
t����8�=�?�%��?�+ES�1�;.hO��ؽTv�1T�'"�ڋ�_��wv�s�6�ꥹa���ݑ��7G� ��ޡN�93N֏�#�	R<Lb�Z	�;���5����ߛ�	�2&#��&�%��H��%�%����PU����-w�<�R9��u�P��&�k⣫��>��Aj��Kk�8�4E.}�t��m"�]�C���e8Y�'Z�L��>HCj`����|������)��`ڂ@ӆGJ4�ܩ.�=��s�w����$ᤅ0��(<�C�k`��ss5$~#Υ��O@U2�]�� �Uҏ�uP?z�ptN��Ⱦ, Kh�R�@�.�%$W_E�9��Q��s��]X�h�"K�C���J>ā�������c�������ԃfz�]��m��v�4�C���e)�Ha��x��{T����(�x1I��~�{D(��ñ5rJ��XhY�^�	��d�Jy�*���H}]��t�|���9E���x����Y��G�4�|��E:�qHC�5G˳��m
�C(9��zj/V];u%�l�Ϩ�
�7��W�K�����9ڎ���f6b�����v$BӼ�ؼ����k�A�м��_����j�P�����8�N|��9���@5b���I�+��X�X�;ta~*�sm���OK�Ӫ�l������0�Wm��u�RX��������v՘>�m��eM�(�=s?D=�z2�� F7?� ��p����$�q�zVn��XG�cЅ`��7�h���Oʴ�ɾJ��X�R���ņ\�0J�>1@��X�#��[���o@�P��_�E����6g!SrMli��F�K��z>�6�)��F���.���ˣ �Q]�����U��w��@���I���̽�)#n�b�ɯ��0�����y�&��AthO�7P�`K䟍� 1K���z~�r�C��A���]�������+�N���Bw|�\����H�!��b)1Wk����L��CMU\`Fz\Yۀ��dǁ�E��^�ҞGx��W
Yl�}
�cى\�b�@u�q��xx���y�kf�[�Kv؎L�y�d���ۓ��]�Hs��U M��s*z·�+���i��9�tGeh(�����p+���E�x�5�OY�_��ԗ��􏴛W�'�3+]�nɘ2er�u9�-�5�����زq�tR)���u���c�,�}�n���^��n�rpG�N�G�����|8��h�V
����
��J�jy�J�/X�$�;�%	)Q�$��%�����9��۟g��gC�!Jj��X����q�ɩx +���}u���+�_�+l�V��;r1��WX��l`z��+�u����4d��8�w�2WH� ���|!����g�xM��t�&ź�N|1�kM>�A�b�Z�zn��[�D�͟������G֣M�T����$R�����'3�{���.�s��������gw`�	���-�Ǧ��U�Y����GNi8#�)J���V�U�6?����Vg_H-4^9��yh}s�&���ю���L�|f���z!<I]g2�7.��2M��)�T�8ʊ�V��'a�����kr8�����:<�{`�w�sy�^�W�6�����������[o5���g�0|�
�>uT�8�y���&����b;/��c���A��ED&[6��ȲgD����"�e�S7����͂7�kqCpp�?�3��l�wy�`"g�$R|��ML��d���g�uWn����/M�<�)��!���`g�r!�'�d�2��̿DI���X�AG�;d%f�'���|�e#�&�fC�ݰ��Ua���b�^��;�ꙫ*�c�n�Xn|��J[|�n�k����x��2e��P�:zÞ~�{�^�	�t�R|�m��"�|��nG�e�x����D�pSz��������w6��V/�L�/�b�Uo�8�r�>�������S���!�����xL��fG�࢒���1��s�nT@�wl��#�_�����R��x(�	vI���j/�Ig7箥��ֈB4�果��
#zr����~xĈ�zB�X�7���P����=Q�R�?��͠r�T��u��	8��[F�0�G?�� T���?C�Ɲm�Б>���n^ߒ�o��3,э�5��|;۩�P5�*�u�s�Ӂ.w(\m�V)�˄�rĳ�azQ	ߓߡ#��(F�J\[�b����va�@T�������od��1�6�ᴎ
A�&�|��\")��"�[���l�g�t��!=��v4��=��CԸ�-w�*�e�;)�����l��g[w3,F",��%58b:#��M����4M̏
�(Y[�&X�(/�O<�74齧��' ���˧�n{�e0#�Qy`#Ȏ������3�k�	�4i_�p1_���v`D\��������GC#J�	kk��%Z�[l�Q��X�a��f�l-��[F��N�u���tj��`���<����`gl�υ����B����.� �:$��R�3��{��=_�(�K5�>�8���q�������6� !�LN�F�i���(���/�W�ep�t����(
6�u�*��F�7�u��ba.�~1�.e+�XR�;�ɂ�R��%x��N��c�7�py���7����Pǆ�!!&�B���fxS�Q��Ϻ�y�������s�;��L��o�
$w�n�.�ų$W��lKm�!B��#��,�٤H5x,�k��.#:?;�g����]<���&Q�C쟌�"M<��7\�(1[b�7cѵ���b�j,[]3��R��K:A��Ou><����Un%�d�Sb.�DW�#��h����$�A��(R�k�s��㎘��̧�X6Dk���%!է�.�F����������Ϣ�O$Z��m�0�b�t,���H����]��D4�1�"������QHշ��_��Z�\�C{H�L��  ���6=׷��B�o%ib�%�zц�o-&��D�f'�&�b"pě�G��f�{��s�o��\�>�P�MiU��k�Z�����!��!s�HP���0Ҽy�9(�ٵ�x�9� ��I"��X�ykmB{A�ɉ��$����=c���F���OȦj���&;\�_ZD@��� �ؾw7F�o�n)��}���JG̕����^L���lB㞪��LU /����D��u���ۥ	��X�!��s�b�,��Z�E��$'4z��!;�C��Y~�?�6b%1�3:��%d��)�FL<��u��o=o�T��H,��nRE�w����~o��i����=�{"��!)U$V���l�ߒ��̌�T�dK	z�牔����4HY%�"�J'�
1`��5֊��`��_9�5 �]��"�>P'��Z6�VW������z���	?�<��N�����:g�s�&W���a�X�����X�ā�����@5�Ow�
'�k�|�h��1Q�l_˚�L�T�i��������H?x+4����0K	��� ��z����'���j*��I$�ۚ�=�p�By}�������!*�e%�U
ѣ.@O��7g������*�B��UV�ߟ����� 
�[�O?�%�����{{Q_�������_��L\���������� s$$[h�J5%)&�D'��y���������2H� k%�>���:b��;&�