XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��A�M�?i��yҹ2� ��j�)}�}X����� mF��%�#po���@�ᛱ�[֐��G'�)r� ju���m`�d�^lX㫂!0�!J�(�'��2�Ft(xI�w�~F��I���ca�!���*y|,i};�S�4dKS	�)��QU
���cY���i��l`E�:�`؁$�UslCw񉖍�����p���hМ1DE�+��2��} �x[��k�=��������s����t�kE���ܞ	X%�ж������	YG�"n���ZZ��.+� 6�t~���M�	�93O �!@��3#34�r�� #FO-�g����Q��i�5��q�ɔ�C&�!�6���񂄰�{�;�I0e �f��x�U*�VF�~kK�"��L/({��K^��u3�;F�{=3jn��mJ�i���B�d  /
/�ߪn8�5�D������_�P���S?\<a��F�`wI�I8昭OD&6W�>���#�~�6�"�s�S�2B��Ӱ��;�4�d�%s?&����%i��B��㱡��&%=
��o��U=Ǽz��N(ͽ���,%oC!}�NXx6��D�|0����F;�$~��UE�6�\y�fI���N`%��Z�g����gu�(�0f�����ɴ�$\^�tFrJ�iZYxr�$q�
%�A�D�{Ӱ�ܤmwS�#_���#%�☆xK��-V�V�HJ��4�PL����&ŐW>7e>� ���3Eh����O���5�vʼC�+$y�9�"XlxVHYEB    dae8    12f0�+G��beݙ*g�"Y�Fn�#�Ȉ����P�9���Hsؾ�T����o����h��F�8B^R��a) )�
M��bƜ�/�f�g�k��|,`��Jg/b�Gv��d���;E���2 �k)F6��+��/��t<����~Eld�EV~1|��pqrcʉ�!
�>�S�D���x���<μ2�ז��VWQ��F+S�d��r��}�s�?/�S�8�^7R�b?�������T�B^g�X�;0���u/_����g�3�_����	�CRI`2U�<*}9y^���*�X�N{�h���N�
����1�*	��È�5�`�2�چb�
pit�o����p����������ƌ� jrj��w�zBg��/�A!U�D�R���.ݸ�\g%.~�Iî ��Mh�����D�lf]�֟�3�>�bA;�v�c���O?�T�.5��K��Q�gS������i=��.v�{�I����p�`��(n��)w��E^&��Zo!"�%��p�wW<Nک~S�{�hC�����"m��bi��V�mcDJ�q����-C޺[��!�`9���n��ɝ��+m��	�mJ5\��C�|O?����|y!��Z��e
ʱ,���:���.͠�Su7�8�i{�����Ζ΍���!���󙝫�J�B�,�(���պ�]��a����>�n��,ΌW)�Q	p�B��HM���(p��K-���A�Bڙ��0
�[
#-�됪$��
C^���e�3d���U��=f���_��9�H�o���Nk�]����&Tn[ِ�������-�~��d���:־����2P����Хm��IUWn���;�3����%��dR0�jy&S&[�l2w9����F�gJa6l�@���㏪C
��hG���P�{�$A+Y��lєc�ƜK�H�/&ф�S�E�r�#�|Svf}+NBΊ"B�x��[�w
ƭ�Y�[_-�|�˩I܀��T�+oc��}��bR��yF���^{(�p���8�0��a����G�����.kƸb��B��~�5��K���1#��Cб~�HF[�C�*J:,[��c,E���%�����^
��"Q}��2��0�N�}ϼ+P���p�ROE2��ۼ�<�> 8�bSW�YcP� o#<� ���o~/��u��M���9g�0�J�ң�	V5�H�9�(��N�I`����M�~���o k8�/��F���[0Ss�jq��vya�T;�eQ���,?=�a���}��F�kM�7G ����W�5@,)~�����W���;2��U��Y�񭁆��l�o�Ѫ���qH��x�>@	rigɅ���A�Vx�Ƙ��lZ)�(1�K�S_�tM�Y�Y>=�������U��vB�QWG-������P1cC��[ERi�n�EZXn)x/ԫP�݈�KQ�9g,7t��u+����b��?�U���(��Hnʀɱ52�R��%��,r���;��xw���C����֗�s��bBb|	G�":Y
�@BZ�O��ƀ��	 �����ŵ;�-f�s*�$��(��{c��h4�(x+V[���'�C�[�¤sy����B���q�j��uyUB�u��t��Є�{�D��������J������ �K�3_�?�&�MZRR7���DkM�f������jp�{#�^@$�_�l��t�}��a���}�_�,�'�O�	�x/��yYU)6EC���%;��0��טk���E�̬�2��M5H5���ɘ	���Ģ�j�����(�ұ�:��MȀE�^J�i�xd�m��Aj��_B��~w����cfqOca��0٫��Q��]:1o��)���D�[D\;�H�������X���#�x,*w^9r%�����I{	��-Q료{L�/��2�Q���_�w�&�ظ8�sꎒ�
&��)Ո�����B���4r�	g/'r/4 y@R�X�-O�bK=��U����ҧ^��vsJ~�`����a�����(	�ؓjO�B���*��l�X�����!*��@�#���5�j�5�cLe6t�2{o�a;��r>^]�n2�(��}���`}���!�8��f�>]�(����߳kG�2h@�nii=.����W>�.��ho/h��(@�r����r�)~΂t?�����<zW ���	��L�@��3]��5il�%���+a.%��KM��<~�*�B���7�M�L}���
�Rr!��o�v��[C����7K�FL���0�>s����b��yo�pUU�<���bs�q#I!�<G���
h�*�fyת�@`c���%��sx��y'840��4����+�ӦQ�N(�`�c�	k'
*��6�>�+v�y9�((Q�M�6q�)�Җ���>h0�=��MU
8�m��.�8�4@/KR�UJU���Z�p�<Qfc�"e�k�d��+��	H�8{F��D�UK�ik0S�����z%��c��,N�Q.M)�	�?Y��Ui=���L�/����= �a.��f�L�Q���2^����އ�R��$�"p�L��GJ
�в�s�2@�V�L/rk|�`O�S.���.gp�BE �����Z��¾}M��@.7$T:گFlA	M�;��~�m�蛝,�J��+����_l�Lo�� m%�7�w��
:tUv4��Z=�����s{��S�0L���G�kĽ��-{�ɧ��$v�Gm�JDB,9H3���ޔ�0���V<�{P�.j,;Ն�l���9~�|����!�����}�qf?��/J��AG��W�\��Ky�Q�Z�EV>�s,��pUL@��o��m��I-�V����v�4\mt�@�Jov�� �o��j�A0�dǭ}�<�J�/��V�<\� �����ܨ��
�i���/�[�JCPx?y<r*��'g	U{����0^�+�$��#�)���6�:Ϛ�VrSb#�FJ�a��]y�B{2BI/�)�;|�b{x�Q0kᙂ@Ah�Iv��R�#4m�$��#�q&���������Ϊ�B�W0)�rW1��Rr�G߻Tȅ���6D8zt�1@RM٨�HA�
(4�:J�-W]¤��ʃDb�]�4_�(9� ����9�n1[9,5,pt3齞;7k�]0s�b���Z�[��ϴ�ո�hЭpI��H�j<?$�-�(o�iV��~G8u�"z�.&�����"���WHȴ�]������ˎ�.��Sc����d�3��	;gM��!�� �Su]E���oۓ{�[��l[h1@��?����"��*����p�Y�p��*�S����JNkJ����Z�ĩ|/�ӿ�����a�<�'��A*�$ڏj^?Ұ��C?<;ಝF�V=�Y�;1���L�u130y�h����5o-�۷���',�3T���-0��.��/�	�[W�o��u����>�R~j�_��:�*اV���h�&�U��Mw4 ���_�����Qu�����Z���u��<0��I�� ��f�q���>."p!�*��+NZ�V2��J����3��jY0� �}	�yr�9�
"��f�#�?I��2����)���)�~L�1��}����_@�i�I����r����+�����Dh�a!�_6|{�0�P�q�i1�}hCvW*>�T��(�c+��,�g���t$��������e3��(�h��Π�Cvr.��e���&T��_ZIXV���n?3I�������S�}����`��@Õ�湧Eٙ���ܒ��/,"�6_�zj��E_K>��ޜ(Ć{`N[��x��؀���5⇣�d@2_1?�L�K<'�x}'i��3@^���&���U��Uc�𼰀#�E/�弿�g%�YK�^��$s,��r(>�<�	R�ղ�M���I�.ے]���xP 7��o�0ee�.�+U�2�	:�#,��'OhC�`��8�p�l������p�[��Ng�GK����:�������};<9�k����LʟP\�*����[{���9ZG�T<�M/��dJ��I,˟����[5ѳa�6l�r�Т'�M&?*��u��_ ��ƈ�(艙l�(e���5a�1���[Ja���[`���.W2�V"gd�b��r������ݭ'y��0Sh���������{.�ұ�^��  ֹ&'a|%�4:`���Q2s�v��"�
kVW���9 �J{i 5Z��"-�`������
9pej/��\T��y�D��{�J���U&�a)��R�nL��6�����bi:��s��Q�>�y����9�ÎZ~�QfdoF�_WP>��l�<��W��"���j(�m B�!�X[�[���A�:����h'���;\R5���*�0|���]���my�z�B�P.wjb\�:�U�i!�yC�JK��)�r���˖��U�u$v3ȏP�ZD<Λ�S�e��&8i���#}Y�N%P~=G%�IRG6�h�Iݹ�l2������x�Is�}!˨�"a��r�Bz��i!�t�c𿣌>6 (�r����A �_�۟����~��Ma �M���!�{����1_벯Ӳ	�5�����A �Qz�/���K�&�&���h���0o�V�}�J�qm���vT��0XPYڜ�
�ti㌂a����Gc��kJ�<�}�,T1��)B.���"G�G��f�\����_�����2�Q�=b�щԊI��
��e�d�������&e{3'�ȃ�s���v̮Tޛ�F�����Rf
mJO ��MAD�