XlxV65EB    fa00    3300L_D�aQ��E��	�J�����=����t��Z6�z��D;#Hgg�z{���hx�X�W9#(��HA��P�H�ú��T�����bMh��L�B�t���֦tNy�����0�čfL`c��_]F��=bO��'�i4��rC4�Aw��}��]�ܬ?X��C��ЎL�܄3(��+Ԫ��	�Nۃ��&_�*�Q�G������}>�R��&9f�;�L�(�T�P�N[V2g᪸&P74R_���XmZ����aZ�����U
�{fM�2L�~;K�vC�� � F5���&�0	DY:���PX���7�%Q!��7�"��)����@7�9�ӌ,�!V�m�#�*����
Q�������+A�$ �!+�C�>[�A-��<��L�z�m��Hs��f^acI���v�X��8�i嶳֙LrJN�McB�IfKbٷ4<��5�<@�#���gh��2�lv	��5�a�[��8��[D^�(u/�!�:���hϘ�YW�4��QEoZV�6A�%��+f��_Ѣ�d
a=��@1N�ZAԃr?G)���s4�y7Ώ*���� ���O�`�|�DsV>U�+���#_i��H�7�a���9Z3���X-�K�n���N�M��h�H���"wD����4Y���ꛡa�}7��I��*�T��߻��<��w��ҝ@j=�{�� ���	���G��1ǵk��{\΃@�R��������E�<��a���*y�+C:�g���ݛ���k�_�7��ĭU�0��q����̶�'���n ��6)��b�i��Koϒ` 9�*�X#������k,�x��1�-�>�����/�Ň�Im������y�d���o-��ߊ�K�.�u}].B�������
���ߟ�b�B�W�98����5�@W��S_��o_��/9)@By�%vU�%��g���A��)�R�^�>� /����;2��À˪�}�Bc� ����p�́p��<0k(��d;��"�V&�	�1���D����h�1u(h  �d�3*ѵ�
х�W�1+�H��$��&OVF�Z<U!�s�z�&�\��H���%�B/ן0�s��O�F����w� C�΢��T�i��8��ܴ�?�r�<�_
R�k�MJ��`�>���n�"�h1�;��y�;��
�:�C�C�Ҥ*
�P\�O ~�
�ҹ�)�&ә��y�?�� R�(Fl*2s��@��#ł�k~���}�v	`��/�������P�ds	'�=��1�H�GP~��6��w̹��B���\�����(��K�*a��/X0$Qᝳ(��e Цp%#Un���Hl mp��`��h�4!��i�v8�9��Z�߳��~ƹ�'{di�W2��!�F��]q�t���(|�����ͬ'(�B��̝""v�%�OHÝ�ٻ�e��r����i� a��ֵ{�ﱻN݀�n��!?8��'����*U�r���OfK����SH�O�R�%Ԟ*��:��-�Zl�"�����꽌{߯�{� G^�tA!	ǽ�hU^�e&�2�iW���r�͵u��7��V�&��Gq�*�(�gk,�O�Z�1�
~��d���֞�idMt�c�,�&d[��e��B��P��d�+��+m��(�i�% &�ӧ�tK����r"}}���+લ��d��ȁ
E$�H+^��Ɏ���-�'[*���Q�����<�Z��X�T\7�QlC��'؜gJ/g�� �8䋖�ۖ#S�\}��C��N"I�R-N����S�#�j�e[H٫4�O��+ ��|��C�/�yN�^�ޛt���.Ɛ������Cꤟ���ں0�* �0��B	Lj���Ad�߿�;d�t����rc`�p@�E��*�˦�GX���eE�Q�6�/���w�텸�͐=d��fE�DfT4
�\��+e�Wv-�u�թ����53���Σ�cK�.��b4\���3-iq%�}1tV��CS%=����%�Wc�!S������.(�k�R"3A�R�YH̷�A5Y܍��\��č4P��:�����������.��H�5ET��Q���Q���q�?���}��f�qK��M�����}F4.���e�)L[`�#o�P3�a��q�t�1�nJ���	T!w��<`����D�@R/�U�)�ڛݦ����)�v�7��!��b?���h�����[V���c�l���,�[vʼi�g���vߣ�e�W��*�'-Z^ g�e=���`D��`���QAnJ�r����f�6x}u}Tw�͜+C10����M򯚪��W��Ȳ\s�IZa�۳���n�\�<�\l�/��@١Hs�h�׾����C#lW+��-�8 �+���c���S�9b�X@V���!�3ho�%Q�5 N�!?��p�x�������9��m������E�Bl�+q�I#A���.���%	����]�nXP�%-x��r���h��)��t��X�cv���S��$�4ꂗc���'��Em�l�Z�n�U����E;t�?��˰.�od�6f��/jS��GjAl̝ΛKf�V~uM*�9>�A_�������%dv}i}~�7G� �:\#�,����sZi�_c��7� ����@#�D� y���0���W�`�~m݆fhb��Aѵ�]�Ke,����B,#��,� ��S�>�x�t cN�o�)xf��䡄4�%�$<́��+uHRq�xw��Y4��8�$�y��&~e妆���#F���(�%=Uը���e��_�j�����%��%=�����'9�ˤv�x!�#D4J0Z6Ʊ�v��J��m���˼]�����\?�z�"�
]Z��#4ڌ8.$�����K�Q8��,�h��v��
���ρ�JЃº���e���H q}���eɢ�;������/o�^��Oq��&^b�@
��H�"�F��P���N7]P��|4�14�;���M�"�:U�d�f����(�\����D܀"�%�c6	bp�Ĉ9�3���t���~J�dI�̉'�"�6�h�Q�l����	�{RƏ�qʧo��ɼ���x��;l�����{���q��^cO��M�����38�ՙ*��G��4�9�Ã��! ��a�������U�>x�0�cn�z��q�QF���v�aw!���<��e9�\�"�f�."XbS�H�����B����l��"
��o����ŸU>O��vD�)O��1YVi)1	��Ј��vL����H��_�O �>��ϼ_;�$(E����.���� Ǧi?r����� 5���/w��N񇙛Cs~��3&R.�HX|�RD�"�J	(?h��Y['᫉�C�[�>X���x���������˷�+@\�����<�t�Ȥ)�M�_܁0�c	g��S��͢+y���H���F���N�_e�gL�	����kH�;?�˩���H����n�x,��u��.ۮ-���D�S�p++�C%�ʬs�]��(';�Ŷ8�bG���5j9�*2|��:A����GVL�O�B�1�?�+��`�Zǋ��l�@�\�؊��6�,AU	�q^��h/������D,�y���2H��+[/`��fbM��<O�g9��1p*���x�8�*J�3N�N�c�Gν#8{��o�H{���b���W��q��j}��m��m�A]�;��ٵ��Ű���#�����aX��@s�+��utG�A
TBזӁ��P�P�ׄn�$��˃�9�zI��ؕle9��'qś���k͞^������j众�80dJy�j!>5��C�U�P���r턥�-t.��~b�A�E�R�kMu%����B$��
x���,�cg�h�%��;�!<�:�Ɂ��'�-b�T�'0b?�Lܖ��ʡ���@�0*zo,������:Z�8�n���68B�'WC�
��4�fIƗE�$XP�#�>��An(�1H@7���f����b�9�9�>u,�I�bɳT�Җ�MC�+�r(/x���N�����-�@ֳԸTCG�xm��j�Œ:��ɱ�Ha#��U�
���Vu�Vw��N����4f��9en$�׉���#��I;�>�b��Z�u�q�v��L �֬vi���!~��mK��b��{v�ݓ��rk����U���d�sK�����g�>�9��G�S��\ҵ����L�X&�v6�a���+aPP�Ǭ�A�'����}�n=�Hgw��Z~s���t����A��I����pBH�/��ŋv��Հ�w"�L	QL��䱕�y���9�.4�x��b�n�$.4Җ�o�O�;��]ꚗ?�cDZDqS>�r��73�Ȱ��$&�5G��/9�zNY��B��v`t�ZJ�I���U� :x_S�1mv�$��Z���Q��k|�?W��BT�w��y�p�s��|XHe��3(p�2���h;����͢xy����ME����!I��r�hR��ӓ؂��=�@;U�f����Eu��r��x��J���w�XJ��^tS��Y?-䧷��F�J/1�o�-5r�\���@�#9˯?`y<&�Ś 9��}(S�Ou4O�ټUf�%ʈ�x(����b�4$U̧-���v.,C��thW�qS�ׯ9�d�DP�<�Te�I��s�T��|��ȶ�fX�L�:_�X�>p#-��kk��;J	=�X����[!@4��"x�r�3UC<b��x��͵m���&�k٧��Av�K�]/��a�"W�i�r��	ҋ�=�3�2�@�9��{/듎�``8�wK�S$~'<k��
�6![9�~�QANC��Rm��u��[<`�S�����|U�S�%5Jl�\L�uח&{�r>��`�B���G�)"�n�'ƃ}Z���!oԇ!1PKi��0����#	E0ēE��g�k�kb6��LXX��d�jG"�`��[����U��Ʈ8Ϛ�C=վ�h�8 F�}9b�������k8�M���|S&O��Y����"�R�3#~��|��i߂ä���F�ik\@�a���'�;�F/SF(`�xO8p����m D�xr1 iSf�֏�+��\���Eb�v���Vȵ񯏖��g6��)�}̣���m��.��^�,m�	|Bft � ��6W��k����63{dMU�:r�)Xq-6&�L�.x��@���j�;<J�N_�]��A~Jm*a��@��9���<N�&�$��4���F���糍�+0)DpӁ�Ԩ�V����+9x��`t�42�A{v�쀍s�S��[��'����O�'*ݳG�>�:���5+��lN�Aok��8�;~ӻIO{8˽@�a�d64F?���tf?ڼ���/���Gx^Gծ�F���Y�U��zG=������V���臠����[� �]3���IdY�(���Da�pU�ղ�:�ܝ��-%�o�˫{W ������,B\p ����t��C6���	8��Y��I5;���R�n��;����J�"f#W�)3b�Kr�3��^��B��b�{�#%[���+�����.��ADR�o��DDO�S��%my��j��K-���c���}���h��ǅ�#�'�v�W�{qj;*�a��
����p.eg��.�#����W�!b���t��Q���?u�qND�Sx���hL�b�_T!պt��O�B���:�X�֘L�|�Sn���hg��2�����h��ϫUFB����Uy�=��|b�v-�Ɋ	�p���cxQC7�djG��oB,��G��d�����SH�W��(�i�$o�0'�2X#��>���UϿH���-�\���Z�M|h����a,��)�"�7�T`Ba
j��#�cJ֧E/�H�8�d��,n��Zf�s�K�:s�yy��K"������o[�f��>�5�m���0蕟@~����+.����3È�����w�퓫�ģ6L���a����Zr*7�.M6n����bx��s�<6���yNS��ӓ%�@��k/����)�)m)�T+=�����a$	�4r���F�]��SY��{6�⟢��G:�\��D�F�w~L^�UY���~{���L
��{��(0��S��������LڛS�7'���H/�.��r��U~c��6��qQ�ܼ.���8��ݘ��Ee։ٶ�=��zǺdq���H��,m��f#b_(��J��L�D�����=E��W��ݻ��p��߷a�|�ΖJL�^L�׊г���N*�}���f����W;j�@x�m�?kx��@�i
ާN;�z�Ƨ��R���{8����߀G��DGO0��N�Է�wp�B��?cH�6����L�^&�Y�e9b��k;�= Zn�5Ѽ({Z��m���j+Qs���Ck�K�����Vœ���J/] i��ً���`���8��>o fٽ_+D��&�64��X��O@"�*殕��#��t��k2�pRۄ�~�vY�����p������-U�����x��z��DH*!��6�Ó=#�;�y�nZn-�K-�<f��V��F�"�l��D9،��e|��Xv�g����x���]I&F�WT2��|y�-���_�D�$�4�2��ϚDY���n��&H��}օ�E�og���|��)�s��G��)�_�]���s��K(Dp.K��bl�f��5�����ӡ�L9+ۆp
-
�Z&�D.�A1��r-���0�h �@i|���NLҺQ"��]�5������S�n�����&˺���v@Հ���`���AR�Ff��>�]�àx�t?��^���'�2 ��6�A��,Z�Z�S�L5DψZmg<\U��h<�ч��u�$��!��|�e�%��	�u�S�����_��qa=�˵Ab	�T �����|���}�h��U��:��s,��p~CQ�a����[�'+?K�E{� cuo#�p�(͵�y;����������'��� ��b��L��!@����vk>�W:B��n\P�#��թҗW�l�����p��+��:�Ôc_&�D���s�_�
�L�J�ԟ�`b���()����2�C�j 4=�*����1�CH�'�+,���|�=T��.i77��.I�����΅�����2�R1Rh ����-�M� �u ��*�޾Ym��Vo�y�8����T�8"}�R����K�T�-V���H����-Tt��9]1���Q�wl�;Z�����6��	9��C`�o�΅or�6Y{�d7�ӛ��O�L �3��.�Ǎ�"R69uh��������,b�9R|ܗ��<")B�T�Lٗ8��v��:��R~�gaE�=���Ӝ��*"���$�(Uk�8�h��J#5㍱� ��}Ō��z�P��Ds[^�lAc��"?.�Y�
V���W�����\�YA87��Դ�����ef��*�������h=sm�DbF��N7o�=F�y�.�f׻i"�Cõ�5\�:O���%(7w���q7H�r����~����I��v���G�{��a�^W��"�Qv�����n�I�!���X\�cif��<\�~6-�g��<#���m৤�/WҮvj��Ҹ����=S*�#�ߜ��fX���(�׎s ��G�P���f��:�6��a�C���M4�7Vq�j_2���{���ǉO�t ܜ���[5�|� Q��m�^?�Z�و	\y%�y��Ѽt��oU���ȫA�.�UE��Ɗ ��;@�Y}��'�L��v��^x��t�ᅞnb_�8��aTg�LH!3#*�N���rc	>��~��I�}ĥeJ�'�i�����B��Y��f���m�m<o�UgI��f�e���~vq�W���O�M�{Fr�4��/e�Co7zZ�逎>��=Q�u���`�'E��t2P�?Ɍ豫16,�{#�_잿1��/�co��P�����K)��:��NO�?��� <�E�Ϡ�E7��-�"p[���*g��I�5��;�=���ݬ��؊aS.PSV�W�יu��t�;N<Ʉ�DǢ�Ԯ������D�׼�2���sYS��[���o�';�c(��4y�X*ǔ�O��jk�L�.oz����ۗ��g+��Q_�c�� 1�O�zI뉏�8j8JBqL>~{�� ����"�q�M����Th,s0+�"��|{��f��z����٤3;#M]���(傠%�Ͳ(��)�G����^g6t�o,d�a�]+Cq�hw�*NAC����FmF*��)�@�� (��Ј��T��2jv��/�}���h��#B�>�,o3x�HPMu��\ڒ�����U�������3��.p:c:�����&��LS�)�B��˿������?f�Ō�B����s�׊d�PK儇6Ƕ'���iHT���������@����ޟ�+i6�^&��s�6����?]���������Ur�nDz~�g����:�)4���^./f�F��x�����:���(��CЌYUo,��,Q[�>5�Ma0�3��c)sI1<h?���%~��Ag2|A�*�01�uӾ|Y��C�n��4��Р�agݖh�3��M��<`>�v�vY���%�;�}��TP�A]����J�&m�m�̸�;0���+P�FǨL8a{�#o�F_�C�_���NHr2K�!Cؔ�k4{��L�"�f�D�&ۡ- �0�5�Ȕ��=��T��#�$<QZZ�s�AY߀��fh�(��u�$�=�8��h�%$ h����ZJ;�}�r����U#��/rQ96��J�|v����o��O$�alo��7$^B�)n��m������K�i]˼Ӿ�2͉��N\��V�cDy�Xr�:%��E�B��ť[��o�u�s
!�%�2�Ҿ���Ƥ�����}�R�1�Wp�ʄ�*٫�Q�Hz�=��<V���zn�κ,�#��)R�-;���٬KP/d�&^#Y}#���i˶����X�;h����Oף&�p�_�r��;0�ɤ�\J.�%�T�I2��V�ܲg��r�bXK��H��Dq�9`�I~���zR$�,��ƺ��QS|�Kѵ��5���8>�h�;%��m�B�<3M�����]�R�� 
� y��c(�Q}��G~�ʀ�	A��dzbÐ@A�q\=m����6BiX
�a��v�a�`}� ����$�%*?m�
���zX߫G���p�fq�N���u�r`v�C�9���崑�q��*�Fէ�w.Bb5���L���*��&�b����IDv�zSm��r�%�hE������h�#՛0�*���_q������?��]����O�����(G�������(��d���II���(jInF;/��Nv
1D��%(0�/��:�K->NM3��)N�����͉`�|,;1�3���v$��3�����H�Kz��)�N@��tu�^��^1����vya��j�R]���Y�����˓�s���m7Z�	�}4�>|o�!�dK��t���l���z�?f�~�"�=_CS�A����ѐ��.�����D��,��g7�%I,~,�5��Jvf'�>��%�Rt�jeU/��i��5��XʻFn�\e�]ܣ�a%_3�@�� �ς��b��b���;t����+��401�y�w(t�0Z*Hl�	,��WSQ�O�$�I��A`�:�GA�Q|�]T�
<��ki˄���72�o����n���^|DHO�k��f=�S��|�}�̔��0>�X]!�!�X�9�3���|w`���6�q�lv`-S��
U;��|F����A���v��Y�c�d��^䁾+aY\)�b�!��g������6<�o��{_dN����Y�l-�J�p�|���k���#���o�#c�����<��t%羰�פ��:��=���~p����"��B�u�:���TC�$6��L@Ǣ�]�o��ڐ�_)r�nc��5�7�Ck�,����G��V)o������u���&�ح��?��R����?��vG}��0� �ٓ�z�1�D�
�l��8�Dt�n���͓v.g�py�J1jR0\��i�]�$��--ٺ�vr��yg�r�H0����Ç���q^��Y:+��x�B���>Ps�Hp�$��폜%R��"��m�����Z�Z���O}ן,����*|t�3���0����qH!br>�`����\�N 7�Ģؼ�]�Jp��KU�:���d�(�vW}��DՉd�t�k��%#r�0dO��LЌ�ҳ;YjI�J�H���� z0�]!_�Js�P��"2���	��.���؍DA������D>�`Y?]�̤a4���$��H�5�{���(���t�/���
�(	�{�t^�>��	j��޹)����%������iV�`]�c�W���[oA��wlB���\��S|�6����!G����Tg��<Rb��1�+].��dw�^�nߌ����a�2����|�w��ԕ,ѯ9��%>?ه�"��R��S���A(�h����`�M��wF'V/ƾ�n�]��6F�3��Nx�\��q�f8;�H�#�����#l'5j�*�H�}	8f��Mi��2�X�f����)�#u�ȉiJD�)��AnϽ�y�^�e���ךq�؛���AM����\s������%C/�"c#���zh��"-#�]��$��(�?(�4�k{��n�@4��[?+/�8��ǉ� }�t���(M�yw��JwA��鄏EH�<���)�xC2�K��\c��A(��W�����/X�(I<�� �6���Lq�Y���虉>���L �`f�(��D���S ���Z��J��v����T���=�]�<sZ�V��������*�LX*����K���!�Ŵ��T���Z�{�4>.�Evo1��L#��=X���O+��g�*v�ی{��d7���� s��9��E���e[Y�����r�B;/��?��`rɾ��-C=l�W�OuQ��Y+i�����ڻj���Ʋ����z�R� Z�̐�t�Efy�.Ź����%ڽ�*Gd-��W���z�ңG��k7;����8���-��a$
�y)h�|Rm�z���滸i�&�d��<Ie?��*Gi����%�Aݦ~�ۿ���x#��
�����̽���X���({<,�/�$��f%����2q�e7���D��D�=~�*5S���6M7(��Y`�����8�	��h.C.�
�ch>��ʄ�pVF�!]ʨ�}TW*�`Vu�0*B�}�$���,b	�i#��8n��Dz�`/��%�P����wr##��b�6�=������j�	]�m�;u�jtu��*�R���[Hi=܌�n���ڍ�!�z�P�*.>ꮯ&��>���x��O���Z��ߩ�%m"�� Y>��/���P@��Ƽ����͹�c9`����}#�1xL#cͭq� s�4z�N�(�q�\�^W7�w�q̘�f����.���&��	��x_
E�,S��L?�R;����^��͡�?x�T[�d��M\!��ؠ��U,:}�.r$y�G���:��ܛ�ɂ�. A؏� �:V银L^%LLe%�<�A|�|X��e�]woc@ �7�|'�"b��ib�6�g���K�;ڳ��ĳ�T�a){D9/��O�]5��ȇ��s��@�,X5�Rt�@����V�Z��v�$��1ځh]\��Ͷ���Яz^��J>3F��ᮦ�)��#ߞTp�� F#��l�'�8��̸5�1��2�;�}X��(�3LSf<�m�. �TK#����������м����*�-J�Ѷ�n��ޅ����V��[�V3�����3@,�1Э��3�P#�������(֑t���NWo@�+j=���X���H�e��/ڴȧ�A�6�V��.��Sx�<;:�z�yX�����'y���t���S\�ɐ|��2���箟�y
7Z
�5 �~��^��_we�,b��x��'rс���C���Fڼ��|S���b���;Xoe�ހ�>�@�����v�#�=D5��l|h��9b���?�r}�'	h�i7����4�r@������@B4��+�
�['a�� `����I��/��K�Z�{#�H�w�T�t���za)
/.~���`�HL$�,����֊
�܏3�)��]�v��Z��XQ�r;yw���)[Ӓ���Z���E��C8��9v<#��MD�:���;Ot����O��S&j�EN_}��~NrOT#A��+X��8�9' S8�}�)��G��P��\�<{�e�q#����ٚbs��L0��V$�r V���}�t2����KH�X!֝u����a�������x��
�J�!� w�	���G�����ӄ�c	�����=��r˪}�[C"-?�\�!M ��6ŋ�sj9�&���suYfH:�hM��q����ߩӲ�u�KJ���O�	Y����ͩP����O?c�e�?4�MY��g̰�6H�l'��9�(ƙ��|�bܔ��� o4)6"�;�tn��OƂ6t�
$��0�҃ �ĲIq��C��o����&e�l�:nM��[��B��Q'~�.�;��:,��?�"5Dū�����H�oo�ו���Ƌ�(8�j�ݼ�1|���s�1��X�6ç\��y�����B���BU�L�4�0�nW�ٳ�[�z���B� ��H��� Čɡ�-�X����������f�^l�\�+t$4�/��qۼ_B�M����?��[�NVy�{C�ƭ(^Kw*E=�����l��K�	�N���[ӭ������0!���D���Y�cv����37d��5T���\�8���yTXlxV65EB    6854    14f0Հo��"�dD:�����"�	c����(�[����u��o�%��-��Ǒ2D����4/�΄Ip�s�*��4w��a�i2�s�ra��W��2�{����F�.�Ja)��8"yȗ���1w�W*��W�ma���)8bl��]�uv"�C��@͕0h�� 6B��;	-�A��E2|���0�e�[�c�y(���j�l���E�
Q��8yK��%�%v>Um�!��: ��6���^4V���5��楘w>((]�ĕ�X�yNT���䖂�2Hg�8)��� n�88�'F&Yy�&�� <�Ŵ>�
�����k&�����G���GHl3�� {�a���5>�.���/˲���w�#�_xs�KM��/�����L^�Y�i�!0��෌������E���g&��v�F��
ivQ�jso�!
���a�_B�c�Z�yS����6�����5Kp�6�w������a&�P��`��:�*��5�T��T�5 E�;�8-߳��QD���Yg���x �Mc#RZj���Ddf18m�~����G��?_�����-�T�kP�^9���M���ek�j̀۱β�<�x�c0:l�{�K�\��Y�h]�R��S�$�C�/[Νĉ@���Cc$�eMob�j�V(�O�G�x����9O��]�_����pك$�(7c�e�]���Ԣ(4�o���d۪j����
'3�}y�I�*nǝ��tt��]:�m��I�n��|����ó�-����g�;$�s[W�q�~ڐ�nJ�I�+߇�)]��	+�'������RY�W*-�=&��X�N�c$�����j ��2OC��d��}�A(�;zbF���]Jp��$<��K���p�A���x<6w�@�\&��y��Q�nW��M9�}{5�uR�T�����S��5����sU@p��oD$�)NX �G����wi����M�yd�D����1�y�2R�it��aa�_q����"�IOm>�H%�m)��8|�i}�Z�rN�j�|��c�}f�R&�ԗ6��꧹���ۦH�Q9Un��>�"�^,���>=�ŊC��Vz)��ar4����wz-D0?���alu*���7(H���C�#�v�R��䰭#���&�&yN��Ͳ^�)���s�`W�k̪�+����/9�(���ʔ��fbcȯ)�`ի���!�&��G�ȓAU*�?���ĉ�}TLw�j8x��X N'1�sF%��}M�?�o1���Zwš^��S��������~Eo�:�c(P���2��<l���DG�l��(��i�6����A�:E9���9�&r�֊�?d�;B�`[�5�xa���0�����>��4�.�U���W��/ػ��
5.7�Ƶ1%	�zJ�7{hz��X�%47*���Fs����&��8��H�MD���_��x�Yk��R�����b��	:VA!�E�M����'#�=Z>�v(V������ <�b��-��H,f)4�0���h~���Ү�00�����!��\y��el��F�0�*��w  "������N(����7�/.�@;�Q�Z���!��9�I2NA�5zC�uU�	���3DTtc��Z蜳��Zp�#�^�̱�v�/�=]'����i0�C�#��uq��H���k�̒��*��%�J���ޚ�sZ`&�x��֐v'�\���P��!̀@�兞��&��_�&aUj�iU��W��_��Q[S꿃�.~����U{J�L��A�Gi�QgD%�`��I��w�,f�3:�Q��G�O4���VLΪ�a�i�;�nC�Lat�Cܐ���4!�_�C�?vV���� ӗ���#�H�����O�X���_Ż��㰁���˾6f���@�6�*��1C��)J�R���N7��Xc��E���3���9�e�_���[V�%-{�r$ta���S#,�j�x=���d<l��[y�4I�����`�:r�	up2K���v\��Y���F�BA�H��8ϭ�Q< .�M��/H-ۛ>��7t�I���U�		7���.3���+|%����9R��l`����F�e���k���3|�\�K�(�x��E�Iv8��V	7>\�e����Xw3hl�`{Ɏ=�]�2��
#"}Xl���S�Ϯ-$=u�5�i�zoE���d�_{��}��
D͊�r�G=�rQ_&��QHk}�������N`�����~[g����U8K�����S�m��@sy�Y��Y;d�v��9:���|�_ҌJ��BJ����+�ΙT%d�#_4z)�(EH�]<vWC��>V�,�Xg��	H��9�ѓI�Vr���O��Y4�WY��st��[u��W ���������J�ng.9y/�f#�X��L4۾�p�gS�Z��� �%_䬂<d��h1�'Y�firOUZ�E��qȷ�������r���>MY�سv���\�hC8��t�́0��^"װćF�Q���u�(�jT�Ks��T����x��X?A��V}~���م�#b��=����]�Eqa�(�v�S�ҩ�iR�M��(�����x��==����r_��Q��epk��3'}�D�x+|ͣ�(A#�x������]w�H��������UR�Y#��xJ��]=-$�@+2���JmJ�E�ݖ7wb�5�ʵ+�X+ݢ����f�a�ݯ����"By���G7S�ӫ��E4����`|3Z��U�lo������d�9��yad��)b�� X��(I����,����l�28�Q 7"��Pf4���}���T\�����{5�]�4d�~Ӆ}���I[��n8��Wp�E�<�ka
�m~���a�w�.p�:Y�Y�S��P7LN�P���;������#��^��6
��R��{��x�/�h�6N����R���(֒/o�E��}�(���G=2�P���Ȱ�g{"���r2�9o�|{F���3^��J����G�B���\���d:����e���M4����"�������y�R��� ��B�e|}C�ؤHk�ȁ�� e���/�3-��J�����XV��Ѯ
�¼Sc���nU�2ܵ�t<p&�M�r,�B�e�o�N�����a>#M��İ�4�;W���1â���$n��Q�K�!L�Rv�\$�@�9I�G��D�0k�T3�@���2�eV�^ [�V��1]��5�W���y��V4;;�<��kd�	���۽�U$~�V[����Gq�Di@!�oB��ʬ���0�^��z(��z�v�Z����+t$�I��ɏ1|����E7�sc	#�]|�[�C5x6RJ��Ո+(kR�Jq^
>=�	 GI�o�rv���y3-��s��ޯO���`�/������JSm�~��IU���?��!��+bF�N��k+HB*R�,�;��I@^�g��� K�7����� H/���.~��?p�5a���E�jNу��OR��,�����������V�'�yHl�4����Nĥ��z&��:g'lL77��ހ�n��]�
:��Ձ��A�C��ʳ8���B�W��#�K=�������nӒE�;���

�Ջn+�*��K���W�'�fs�L�*IVW�-a� �����d��%�N��$�r^���B����2�".\l�7�8Fqq\Ψ��o�{W���")��i�"�2H��hK�Rn�d x%R7C^��*��S� ������hc���e7��60^ش�#�F�����O�-�vLĶ̵{�4{�hbt+�) ō�Ȫ�/�����D�
�ţ2�~�e� ��H�|@����_?�h ��0E�VaG+������q?3���H<,V��X��嵘���f�����a�t��X��
�J*��e��1�	Q��ѬZ�p�j�d#�X�J�:�/<f�r�h(n����U�E�b�Yo �����$Gy�������ށf��vE�tb��싥{��_��u�+E��V]Q���( �0�;�[#P��Ę��PGT%�\$;�E���K��G�� r^�KA�t����qƛ��
��,�=#I_�+�>�~�����&���ؠz��Z�m~�d��o2&H8bK w���ӿ��B��&���≵��ȩʃ�����t!�ԛm�����}�v+�zƱ�� �dCbh����R�5��P_�Q��׿�A����l����rF��g'U��� �~�2��w˳��u;��p��	~y?�I��*2���F��p�4�=��HYk�ƛ(���<a3��Lq��n@�>
��uI�6��`�.YĒKFw�\�ϴ!���u(��U�h��S��xJ���x��\py�HH��O&3A�0cd߳��+�+ �����,���̮�*9�����L�¥v>�̞V��6!�|�)�@���c�Fw��?�yVDg�G�k\��:w����G�=�	5��T�"S=���a�6>���O��wl��ز�n彔3����Db��������߅�״����w�AAN��Z�fQ����h�Ef��ܧF��:K ܖ�\w=S������J��VߙƗ�� �׿v~��+��*�b�v�Y4��4Yo|tz{�F�C�u��<0	Cc�A^6X\�s�Y����ji����HT�4�'�����	 !���=<���>Q����woM;+Z��Z�^�R�w�'�ͻ��+6K�G���FMv�Ef�ʚon6Δǿ����?�:�n?��*8+�'ښ}��#?�a�ܡz�JA���&��T��g��'�Pv=����ҧ��f��"����A�:�@&,Uj���-.O�>�:,�˟f¿?�ᾙ'^����7Eb[�_�[�-�ĸyEϙ�m4����!	�m�"��
�>9?C[p��i��14�-�W�~eG�l�u1PS�t��1���֣x�8�E��Ľ{C�a�l���R �Z�W��.�g	�2��� �{>b�_�奎�⿂7�ή��}�5Cc$AFs�4>O��
�
q��,�rKդ�������'<��3��5��pb��E��;<�ȿ*���(r��'A@�e�O��$�<�����W�!��>$�^
��IZ�0����s�[�8I�Y'0"�T.+B@;������8�q[��j��@�f��v��Do�ZA�Q��nU-�,ޮ"s.M��}�\��c9P8�*
�a��ɧi]W�k	e������
/_
|�v}CA������{�a��_~���O�gI%|����:��}��p��G,�	9�0A������x��<������On3o�@