XlxV65EB    6b34    1350)Cs|�x/�L7�u4OW�����ָ��,s�D��S=��*s2���|��ޏ�������[�8����@���uΦ8ޏ��;�nAM�%W�`���ԩ0h��%N7���f'd�����Ő���%@\�<�1�H������E��>U2yb�%�qT�5�%�����<���S�n�z:�,��G�q��#�r]/ӣ��3���� S�����`�����̻�ݍω����;���;t��o6"�v �+%������x��yM�f5\���Pk̃: ��Ƌ�e�̷*m-a"���m�
�67����O��[�GaaB5q��K��H�+�[��g"��ǔ����!k��Iؕ�u��O�ۨ�������d�n��l֭���1��QՒq�E��w� �Ƹaa�	h0߸�ڮ{�(��"��Z(�������q�1��J�/���fյ���W��༹�-׌gP��bH/<J��bL�-�����̻br�t�忶�8�A��=�^�3Pù�0��e[����֘l~O��s�6&2�(���]��.��p�<�49$�F���Ư�E �`�C��+��t�mܹ��wG^��*o�NPh��N��SzU��(!�~�*�H����֕WB6�~q����!r�3�C�~�&Us�b���q��Tu'N���#FL�;
��_W����-y�B�Q����hP��l����7�����'�z�\İ4T|�6��ic]�Ѿ�|n�V��,��!n-�W�&�r	rÛ��N2c�F�nK�I����/��F
�(#�偁x�(v����~ʽ,)2F�� Tt����Y�����["��8����aak�}��-�PA���Q��"�z�@c����/w*�_����R4����+v;KK�L���sl���3�q�MU�{�-�p��$f�;N��5���KZ��I���7<f������I}��~I��"�=uZ�*Ht�;>���2�m�m����)@)���kE-��S�g:���Lc��*�W�����i8�����nd/��ve#Y��������l �������Jf���<�>S����r����lנ�}P�-	
[������/����� ^�H�l���5��~��r�:��h��~���bG]JB���WE<�����?�J��µk{��`�9_F�Z7h�Hv�Ӽ�Js���g���m���!��\u��g��u�AP`��8��0�d�1�\�B�~P��9e�w(1oܦ ���]��O�#�V�b�}wT)}%m���P� 5�}�Pɶs��T�5�;�z��Bp@�:uG�;�4TK��ɣ�����[u�VX�7��DJE����rL���٥T륿�/���$����b�u.��$s���4�Sa��?xKE{y?%g9l�u������?�e���tļl,&w:A���TTw��K�S(��-��7�N^���FIr8��w�O�����S��tG�����7h�X�j�;#�mA��x��K%������JĮTkb�X�NU��|�8/Z�F2�����muL/D%tl[�@���.T�1W��ZlY AZ�4�x;���\�0���s`�o��e"���V��6b�6%��NE��DU7vf"����V���%&�r�"Ӵ�ϟ��@4��\գlDz���f͹��@������;	�Hm������¾u�@�8 ��]����$�F٭a��9S��פT����� Qo+������Zx�����	����5�R�i܈�t�#YN
Emd�D������^��`�=,�1;gf� �u�>w�2wa{<�p��<�xT���Ġ���I�{7��&�2�Đ�n
�Iy_�+�����\98	����mS�T��s�%���r�㯟�΢[�ԨB��T[&�-dK��s��7�g�Z���i��G$� �����`R�p�c�s�I��]�ZבI�z�Bi�ٺ��!eծĈ���^�"�^��;�Ue��l)�S�|��&+8����:4u��Ky�t�p}���Sùt�ݛ#_jRY�2����Y�8���%[�c�`l�G�m��.ƒMG<Ȋ���
��$�����=P�s�!߱jtu��>�$�����ks���6}NY�[_��C�2���G��%�����Pp�゚�[�pc��E��,@�)>�_���vpW�f�ژ,;̉���xWGA0�ì���\D,L0��
�rD��a���}�E�i�a�8�����R"vH�}#)��s̈́�u�-�O�RN���>��J2�.1:?�ݛi�Q���E7��՘0	�P���U��O��Up�W��q2�?]oa2
3p׭��jyk��u�k�k	�q�Q�ϒ�ƀ���	R�6OȤ�:,kJ.��}X�@:�nTQU^f�8��^�;�|���������'��ͽ��j��K9��@)��jl������������!D4�����DJ�D��*�X�Nˤ����A�#=�?pz_",䣌��<e)Ɏ�`Dr��p��'����XJM7]�&m�gU,��YA���Oo-+(���%��\����(eq{������Ə�	�`�T�L��~���"H`l:'��}P�Ѫ�Ձ>�P��7�*Γ�E9T�(8>�#�7����)OG]�� 7g{��L(�8��v�{BH���S��6vl�������{�1���E��fIq�a�(B ��3�+
-N^���N?]	~��(�����#�d��>�����o↏</}M&n[���8JV�heKD�!����<�:�m���EQ���/�}0�A`�����Q(��#����>>�vvL�E����%�X����NH�{'%�<����r��T`l04�>-��SS}�+�?ԝ��&-3)�҃#�.�<�`ڝ1$6�ă�@'����`be�F���_��%"��%L�c���Ǔ��g���jܢ���k�Ѣ�O/M����M���,��v�W�RC̯���J�>΍0߾�S��'� �?���f�5��+J��?_��F4w�`�CgF"�Q�aGp�^>2�tN�z��_�7e�P��&t��0D�X��Z4�����$'��Q��#�p�bCz'٦�K}��\��s�oHS�-���9SG��#��AjR��<����Uɠ�|5aVe��e��eWa3�V}�L��l���m�1��K�W�"W��NL�g	3��ξ�읩�M� Z�3\���[���e��3��"l�:��~B�����z6��9���Q��F������i!�[�sc�G�a�}�&iDɅ,��XЎ�?ҪG��Jri��L����ރ�w�[�;�q�F���H��XK�)r�'z((�V�������k#oz�e.4zs;kG�7��U���c���u�F��	KI6nU�#�h�G�n����9dL�8�#W�u$gB/O�����Ipm�Ԋ�A�,�����q|������
5!Z����]p����]҆9!S�M4�4�.��ch40��7��ெvS��ؼ��i"�h:JL���;8�nmѢ2Հr���{���Zנr���������2g�M���>KOU6B�A�ieC��R;��ݖ�t�)���Dx��hy�
�s��󵜲S �=�>h����}o����3���Xj��%��.�=�?w�}��X'Y�=������no[��lO���5 �>��,P�oI%�H��?�E]@,M?�$�ǚ�)펥�i�ix�e��vo2�R�ݗ.�4�L�*�0����3~9���G�(z�׺^��j���Da������zp�LmȷkS�
XH]<�޼���f|��^��%�D���k./� �is�@Z�
D �U�la��k^�����W�&�4�}��k"��(e�׃�ޯ������k� cv�`�ǤX�]Ԙ~@7�٣F��J4�����_AxXw���U�F�lܯ0 P�s.��xU72��/*�j��-us%�fa�p�X!x�̫k��F� !��B\���z��Z���/m$����GHH�<�-���sX�y~�h�G���L��ugU8��A`Je�!(.�/�.�sʃ�ǂ�ѩ�x/���Z ��
~'~5%8�)�{yr���:ݹݗW{���Y��&~���&�$#�g���Y1\���|������4�*=��un�l��E��K��c,Ɣف6Ere:Z@� ��dgSt���\	��B ���fl���ge�$7r�����3�f�^��Ɍ���eu�l&"
(`^�Z����_H�ыw��������hr�m��� ��t̖&�j�O[�ϻ�g;㶁8��[�c�݌00��ȴe�����qƆ�Ͳyg��u;�bX����uLŠ�s>���G�fʚ�l~��V��z��3��d�>w�b�_u���f_f]�F��iD�b���gN���,�{V��s/�`��HN0T�C�E��肗�ax�]���Ǜ����������F8
J�DX U_���!�"��:�j�imgLR���g+ �ϗgF=�F&������O
2 d¤?w�?��ȼ��P	C*��&˶��c�k�3�O��o>���7�%Jd��w�������,�؀,x���Q٢���W5�:(�Jw�)y�#r>B��0*?}j�*nR#2Der���7��U;��O~�v�EՄ�hdU�8eou7o���$o�qz��oT˜��v�:U�%4�1BgN{t�:m����]<N���u;kѲ�L�����6�w� P��Mr�
�����H
y�(J�2r#�5V�sLh���9�_������ް�t>����S*_Iʐ��%~��Ԏ�ڦś