XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���%��*�}��-d�L��7n�o�}'8"s@�c)'�;Ў�/�ԟ|#H���܊� ���\����G0���� G[*ˁ/�D��`��h�������JX[7s���e�q< �^�a�	vD7�͸̴�&���w(��s��+Im5l̎x��@����5�Hv���|>Fe�^�� Xv��Md[�HW:#��@�p�����=���0Ij�)D_�|��F���;vޡi+��mm�N;e�"S�$�6�Q#�x��ox�ω�r�hf.��򶴶�~�]Җ[���P��}<=���������L���Ƅ��c��<-R�&�%�c#^���2�.����RU|1&��
'F�/�Q��.9M�|�l|R�O�]I������%G� {W,8�Z@�����?��{s�SM2-�cxf+K������R��6�J���l�����@hv'{���ck~m���?����m�r!��]+��z_�Ӳ�a �����Z_7�;�Q�dm3m�Q�c�����M)��IR2��iT�s���d-G0_o��|1���?��-,�-y�-����%���bLM��L�m�Ĺ�]��{Sַ��u���!�z��|�p\i�=�4]p;?}�Ii��p!���CԄ����%���Iν����kA�V��'VA=�h.0ݜ2kB�I���o�r����C;�<�#����� �7�@����K�I�c�H#ħ�<��I$�h�~8;�iߵ�~L�XlxVHYEB    80a9    1880�J_��@+4�Z��I)��Af�K��b�xd�T��f�W�OL�@0�F]T������@Oʫפy�)�v9��i����G�YF���+ uQ��Za�'�s��6;�)��kbF���{�&��[�C�Rd�3���M���-d���g�q1/�z���)Ah_���h���Y�����y(������ű)R_���d���.����8^��ߗ])cj�aRc�L��J�Ui���@��-1{���ѨN�W0�<Ҿ��O��/ �+���M�!�g��OC�����m�-F���V�> x	�1�a;G����;���7sޙ*k&��3��rpB
O)�vۄ8���C����h���ȱuu?W��}�$g8�<Cз�A�rg�)Y������/�S 0-(���T��xh� %nh��h��m��S�[�%7dD<A�%ܶ���*$l���=̎X)(a���F0E
�ps%�"���]
[��3P[o�z���*q?1�UO�z@�����h�W���y!�L��`�Gs�E:n��-;��c��b�ؑ*CU�\���BA�1259�K�&�m^�u@��]
�؂#�?WRk�,�؈��q�"��z�;6P�,گW8�xg�	�#2�w۷�۴���} �ze|׺p����{�ش����$��:�Q�H��yל���)7<a�i�oi@"����X���m�YX���ٯ�yBl^/Y�p��q�����{��9�%�#���)��L$�BM�{n��x�����%�\imXx��{���=��@7:�<L����38�V/%.3��U�ٛ�i�<L��͕���?v>\���)"k���Z�۬���-Hx�O��^�K�@�	�D���I�`"ۆ�d#��?�M��W;>4ߐ�B D"{�e�S��A�]��3�+�v܈�'UZ�nM]4���J�����M��1��{����]���w�,:����:r�7�$�/��
p��!�50.rH0^<0,t�UO���z���p���Y��[0|�D�y�j�3*��C}�	�*�7���^��TS-\��Y$�n8�������7i4Yld�o�~;{<�C�inc��}�ӣw�i�sx^����G�Z=VI��s�T��A�Z�ps�qb���U}Ǩ�|��L���G����G>��)�eG��2�am?�Z��z=�pX	\CU�4���{�q�rǦr���������X����K^yP��9}!��u�����P��BPjU��<��m�G`��![h������3���`�&��M`Q���F_�Z
�c�m^�1u�P^�c�Фn�j��^��n�A���(�1g��&3\��i_�K��M�
h��q'�V��K���P}��U��	4s ٝ�Aヮ��٬E�I۾�П��+�+U��K��cf~./.�r�A�eʒ���<��
�D��������Hͮ��>�Ƨ����c����ؿ�8�9|�,��,�����p��e�JM��e���i[���-e�R��z���|�^
�.;*`��|۸T>p[X*d���2�[���7.������������?�y/Ux�U����4p�ss':Q�@�x6!ۺO�T�b	�*a��l<~�a� ��e�F�[I�,1H懻�Rv�f4����tǎ�H�i1��~��ߪ����{I)Ⱦ�}H�(T��Q�!P`5��1�K��cK�VDG^>i���z ;)Ń���v�_$��.#mM˘H'1n�x�{~�?�<�Kځ��8�m�"���UM�����r6��")����YSi%�ب<g0�Q��l�皉r:�
�a?���zbk<`���fv���h1���~\���fbca��~��Ȋ�%f���"e��>��~���q��N�x��\�6��޸���Oa��a�gP�f4{R���]�i/r��i�H��V>�w�g�o�W�&ݟ[f��� ��=�o���	[z�`V���MW+���e����(�tyʷ�#���;����)LL���v��f5,b߈x���r��-�Մ\w�����9F�6 �E��J�����!D��
jj�S�O���va�L:�)A���[��<$��&�\n��b����XC������_���G���z ��T��]���)P9�D9~��� ���!���(s?�5L�J��*�a��v
w�V�v�qeF���~�+���6�Z^�H_��3'Z<��#�2z\&2�XlB�¸GZ�:�5�T�.߳�7�1�q+��~�D�1i7��չ���0�&�e0_6.�!������A���P�+I�Zֿ ,��/��A�,���"1A`]M�L�^?`�I���I$�W��%v����(t˨pg�$��!YA�W�#�RsP`:9�+�s��{,�2����P?�_3�.��F(k��y�g�:�Rv�j����U�B�۰����������!�޳�.=��*L��4��ͣ�qx�ғ�lD�6�e�^=�����i�Fz_� :�Q�Kh��3'�}�?���hHv�h�eb��]�g�]%]�6V������C�iK�z �=��7t=� �G��M�D�Km�+t���zx�p b�����������%h�.Cw�d�N�t����6�(���bM�S���^pM+�C�Эi�/�`�#�G��蔙�^*��o/D��a�1��RADM���4/z*F��!��R�X*��������dЅ�����O{��X��b�z����G.�_	����3 QR�ǭjN���Եy��@z{7��p�PY�s �+��;9��tv�H���Vr|?�[��M2�⺊�};�vP��x43=�@����=�~M�չN����u�=E�z�Q2�$�
��v�A�EZ������tZ�UV�<�w��[�)�K��i�i�!��p�*a�T��fRЄA0��:��+C,ӗ5�H\uj����f�b%9KZ����]�`[��i*w��.x��\��`l��QSacO�����l��܈�����*��&F�jH@��[�jB#C���/�)�b|��N�	�WT�د@�)^��0�}~���59��� Kװ٧��r�$yA�9C��J�N�mpIH$C��J�~���nO�<�������	�L���=l��wL�*Ϋ��. �����]����v����۸ѭʚj��5�k�9�4��p&�Q/`܏M="�[�����mTIv־�u6����e�cBz�b*b��Lé��af�����T����J�O�e?7��1%$�MF%�f�Y�u���v��l�I�&@���B��v'
�ʢL�~�;�U�/I��b����H9�Q�ag3��M�:���f��+}mnsm��g�}]h8;��R�B̥n6=;eFy���ٖ]H��P��𝆙t?	�yň�C߮_ٽ%m�?��r�&U��zO���>;L�����W3F�5O�^�O���'�&��3X�$��Z$����M��ck�@�`V���6Ŏ��7��sa��ȴ�qAra�l��e]���J�T�9�.����B���M8�ٛ������֮�丒mb
j���Ӈ�ƭ�]���u��@(;���f6GZl�U^�s�g=z�F8�&�2e��Eg*��7���/���+NYg�u�hዙqmQ	�6%V	�[�PHl�x��ή�	��>$��fW�ŭ��\������7m�%`V��G��b�\]:p�ҽ7�� ����+rx���^gY_�.��&dЈ��|�w���/��o��#f`�d��B�o�4G �%D�̕�P/OpKv�l���)
8V�"���`HhD5P�͕��-u�RQ�=Y��;�}�Q��������b��
S����/���G�qg���Ç���z��7��^3�\��Κ��L�����#M������Ŀ��5 M3�a'�笠9��y^M���о�o$z�\�VA���^�������Z&�C�-�A��N���>u���&}A���9ļ�鋍�lX�J{�MH|�˹Xw���� ̽���?gt�������m�<XM0~�#&�z=%W�	��5n:�p%^����g�b���k��A�O��H�7>��7��x �����5n��P�ɨ31Y�DpnJ�ŕ���-^�X*k>��^y|��;o�!5�p���C{Ul�VA3�>�l ��/h��J����ck�e�_���Hl�4㕟�3���Lī�f����r�J����H�?�S��Dw'{��]��TQ�bQ�DP��j�uE��� �X`4���<��x���Jg�S38����ݵiܠ��ţ�j����t�`�P����8�=�����=8B�TID���L�״L�N��c4=I�Q�$E��=����hqs�����T#F��t��+���,>@��(�D�3$��G:��������n�]:s����N� �G@?���Ax��n���T��h���G�W�I,K�l{�H�S)��ǰ�)!qޣ���]���ȡ�j=cE�U�ǣ�̿��7��DW�Ri���ɷR�Q�a\Ѝ�a1�D��JO���_%�|q�� Q�7�N�?�Tc�R�>��-4��|#�]�n��n��S8D9M#fDr�}�0_ν=P���Wh� a2%�P]�)���-�L�c-��)G�Ч�3:B��ܐSP�/C{M���[Q	=�L�|��&4���$#`��WP�N�G���3�M����#��Q{R��r�N��|u}����6|�a'�0�\��f�}��+��?Ip�Jz�������P��z����1U)��2O %'�����-?�WB�=����N�_лg�p;�3Y|�ѷy�Vj��x%�n��'�U�^V�VA�����yǷ}%O�b�k�H-�����<��K�$n�m�1NF+�����yav�S���'V-i.�:���	�%�&K�غ�������f�����\	*� ������U舮ڵ�_a�L�~�֐ja׮��:��ikO���r�Y�:���S�}�;�p�%��f�^ ��.1�ET`�z�$	�<�f��߹'�u���$H���E����	��zʊ�5��($��xi�iQ&���ˉ%>n�!ē���u�gu���~7�d؝�����,���W|��N,eK�q�s�~e�0;&2֝#�să� �ۄn�Pu����7��՘b��p:;��9�c0�{���_�C��\��C���E	qhq
Gd�,��7y��n���	4׋��R�)�_M=1����<R�N���-flR����U��Bc����INF.�NUE��5zI��ħ,'79VHGx�7�7�>���J��5{ܗ8��Im�v�I���-
��0<3�w�A�N%)�Eg@�\�_0��4��-�q�w4�@�ش�����q\/�3��$��� ��x��7�j�o��׬F�=���1�%}�����5���O)�֙���
'�a�3B�T�,�1g�0�_̦��A;����Rq��N�8+1��B�����V�\�F=���Bx2*��!�KXi��B�-���d�`P���.�g�XS߯i�ج��(9�B$�K�$<��� �\���1]uxݴ1�J'+���4��_O� 2磻V����Ǚ4�;���=TR
�'Ɏ�����X���/��:h�ƌ�'^7�sZ��T;��[����T^�.���E�{ᯧ��]^��X+��S$iD���BA���_m�"ly4i�-~@�)��@�r��;����	Ev��1�
�
޺4�?֖̗*�t;�[A^�A5��\*z��/�����ljn���Ν���� ��kD��O/�h��Y_�i/�5$��R V�BNyJ��V)���2�f�19o�B��"g�>�[iT�3NI��0�˻�e�ZIO����]g/�%=6B����(��l��r�4�X��D:�Ӧ���"{���p�:+Y�ݛ�J&�Z�K+�J��XW{Xy:���t��Uю5	��*�`�S�����b��LM���9�d���dEt@ܸ{��Pp:J�~�֙-�/�<������5-��l�y��g����Ԭu�GS�-���vC��8퇪4o�W�4�$.w�d�H�m��쇥U6�?vH>���4�H덭YiѴZׇ��٪πd���D��������"ﱳnd}�W�