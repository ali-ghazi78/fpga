XlxV65EB    5236    1310Jd�8�(��d?��64�b�5a֋�?�h��I�Q� �}����+	��x�Z���y���zw�V��|�*�Y��������rh�Ӫ�<����N�b��VOn�����:�bC�d������:_?[y'�P1QT��`F�����ܤ��to�@$:��Ъ27Kw�dͫ�[�+�jt �0�4����Vg�y�y_�#���j�(G߭Lj�s� Ω�����m���oLJq6���5.7�;;./ȡ/���l��ӽ�|�9��}��������R��$�kx.TZ}�>,L��ud!�2/?�x��-u�d��N�$sO�'E!.5zS��y-�ѵIz�M�۠�^uTn����d�)����w��2#�m"��a�L�&�`N��=9���M����1�y���!:jR���)L����ං΋�B �ZRa�SI1}鐤��w��f�}�x�$�Mw�w���>�N{a"C��"�u8D��>q7\�Sߧ1���������8.�b��"�L.�-i8�Hx�,ܸ��짊���F?�Нo��mk#"�l���g̙��O�p� ����3� }r	6��M�3
'	���f��$4��ΡQo.���x���ݕ�N�N�9�L ��w_�c���u��n+W��|JԿ���!���� 6���V��.���8�D��Ca� ��"]@��ܓ��r��f,/��,hI4-��n{S�>�MJ,	s�)b����PQ��1P�B�Y���y�H��A���.l;=]�rp�W%j
h���I��?= ?%��E�b�8�;����I;��t5m�ki5Rs�Ļ�
�̦���`���C���>�MR���x*m���!����]ƾa�,���]}�"�uT��Oq.�nG��%�G*��>߫)$�>�Ф�3�A���"���vQ�F�D����p'!���z���
�Or�rǑ�ґ�� +I ǳ)�my�\A������uҰ�g�3l˄�EK�yv�+O�����!P�5N�I4�/.��r���?��m�>r�tU���L����"�v�O����F�P>F8!���d|x�5�r��,m�B�ߘ�o̢�-��W�X��K��EJ1�2���M0賃� ����3��׶�y!�:J����ۢ>5���I��Q���|�Ǜw[��݋���];~��S��FC�7)]�<�h1a,oȍ���` �-�޾7xԎ��iR���Hc"95���f����F�K��ÌB���s���Z��@2<��&޽0���3���c4�} \Ni�6�H˔V��>F��&���j��/ou���V=�z=�m�EV��<�0z[P���P���l�ՙ8����%�7���d~�����8�`��c-�mn	���7��$,�%�<QS��a���!�h@�z��k
��5Ln�9�*ci���_��.F�Wr:��}4�
���Ł����3w���e��u��3n��|g��8m����+�Rá?Y��R�D��+��+6B�tt�b��l��-�5���-�@��ūcR��&6X���Nqm��Y�y΃n�#��R4��:�:y�=<z���6���#�U1�'rgP�C�3���a:�=M��؅�|�����k���N� ¨��PZvy U2��	5��ay٤;p��n��SgX-�\צ�����j4ܿ�Η������9s3�j$4wR�o�4.�1�-`�8D�k�@�4�*�{��S�钬�2O#��CUF�􌀔r�Ǔ¹<u�Y��}r��`��*Uo��1ey����+{�<\�������on)��D�#��&O6e��վ憊�Ԯ��hv���8���t�	%���v��38�@(�C�t|��Skl�~U/�9���J���͏���Mƣ֋��q��IלE~��&�o��):)��ZT�L�R��8�؁�c�%�c�GK��x9s�Q@"PP9�xp��ϏY�ĸx`�ęNVz*7�󸫴��t�����9�\�0خ�\^/�(��t����h6��{����ǈ�~P!��Ih���n��Bpe�O	�b�_Xo��!�ө��R������b7k�n�A�8�u�&�Z���aY �Y�Y�@�)��dAV�5�E�F '��Q)&���yBh8?]��Z�__ f�1�o&�fD[�#t6kW6hF�S@A������#7����ʜY�nm���O�7^���+#�Fg�מA�p�����
�"=�R�LUE��*l�Ҝ�{*��ΡHe����Y�� �9{�7�r�'<�c1��&�kVl�aQ��C��ۑ�BXG�*�<ſݙ��6�t
4FKft�}��Zfu��Yy&�m�  �zU��$�2s��Uz������*�0\ּ�\������5	a�[%��>��%���_�{�Gc����x*��i�Ѻ���K�D�� l�O�D��]�r�ܞiޛ�7������]���l�2�@�N�5KM���"���1�����N�Ԟ�y��5u��d�X���X~	�z�D9p�ǉ��}`�pb�
1�j�،�/H}.���@��E��M��ʰ�����p�p+���}�⇛��4i�� ?��n"��K����(S>�(�\�y���us>�{p̽B7h�
��K���'Z�Ԉ��zd�3H�NhB�H�n��n�@���9��{-��ܢ�~t��/yp}w��3)��AI��}�H� u�������S�#6|�y���c�ܢ�g�uԎC��Yl�"��?�����f��B�GS�:�J�K���j���`R�SD8��@�����.�iCnC�8��������{�T!!��F�sV�г �p>l8�73 �,�G�3z�r����w��Yj�[{
�N��r�-�����uP����3X�g+^U��bL� �vHɰ�d$;>�`A?*V�W��W(�D�i�m��C��%3��eP�|����p�;~�h����b�ݛ�l�b��'��)���zI��?u�RZPw>�>��l�h=� J
c�=��z3�F��n�۠k�5 N��P o��A9�Ch/h�I51�>@}�s�B!����o�Yb�=���җ��^�1ڀ��[�G�9����9���l4(�@$?�@�M���긛i���4ȧ���7ɗE�@�ě��������6-��5xU���~;!{���^"��*%�� �~�vAH�����4q��5��ذ "�d��& iE�@�4}�`"�z�}�����q���lS��f������X�kM���,�x�E�{�L��2z�S�ӭ
4�#�����v��f�GM��Sr���'�6G��~]�2�Yꁛ��:���gؽ^u*F��in1�hހJ7��n��$GK���\� �B��I�����Mw����;�}PJ���d����c{�s؛��4\�M��	�At	I�$����Wm���D�㏥���a�/�(}[����`#�oJ �\Cjq�liO��R�(U�%+� D&���)��E��X} �?C�K.�k�������ƪ��	�D���5�����#Ղ��2�g$z��'
ib#Ը��,.5C�vZ����uk&^LU�-��>8�ڨa:���>���+;Y(WB���%j�W�@)Z�$�O<3
��}nXG0��& ���k�$���ƻRb����!q�쑐TT���:Q#�~(@�`��+Z�TL`;a^G��2!Q򪏗���K�|]	�V�н���M#��D��*|�ei�L/��R���H���/�S%Sq.��5nM虈�=�5�r����98m�}(�����h`'D��X��7A�s���%}�-�>�	u(��?�T�!۠Z�ju�	BU\al',�ӏ�*8�'��F`�2<[�5���$��	�d;�%>�X������-YC3�~��8�7E��UO��pvn\f�Y���`&3n.<6�� �\���������>ا�U�@�~��Z5�`P'��PR����P��v���L��D����"Az� z�5��_qƋ����t�±&c�?DM!եkvlS��Q,��H>����*���	�����!�ҽPp=��Yѻ�����n�ZK�]�_SS��LjF+a�������a��H�]A� �k��K������0Ł��Bw3P^�����`�p��Y��n���怑'�H͉��S���`�2U��)�w�T&Jh=����V�x��}n���-�;��_DL�@�>����Ҥ�W�lLK���B�b�#�|�/S	d@�s�dw��`8)rԼ�m�c�̌�C읰��į�2�퍿x�J� ��֧��<�Mc\4帒E�F��gݑ����r�)���.R�Lj�~��Q��m���7ṳ=�0�
��l�4(����WwQ�¡�`Zێ}_�mv;���)���'=L�{έ�N�0=���ׯ�c��W�]��������}e��խ�x*�%cw$\��R�E� N�s���|��Ub:P%�)S ]|kt��O½0n�c�q�e��H�۵����.���;�����i�B�#��hvxDo�wf����M-���0t"�t���}i��N����@�&�4Jy^��c��4_W@�n��Y��c�W����ex�#y"	t�~1<��!�q��"P��}�/�
$V@4s�[���O;v�9�9�"D�W�l�y+%Q%��ffpYEס�+/b�� F�O�a��g�UlQ� �+Xw{�y"�iB��oA�x��О:�͝z���v��xg�n�=B�lE��i:��>�~�Z���ԥ8�,�Is�򉾨�Τ�#�����#	M�LL�zϜ�;�da�`�"cZiJ