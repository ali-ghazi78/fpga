XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����#�8�w��P�H$����伫q<��|D�0��<��QD.ڳ��A~����AO,��Pص��V2��	�=�N*?��U$9���,ע�利�*K�ɞ(*޹Й�J���;Q���m-��ST9n��G�����ߓ�9l�i���<S�	_�z���YG���){s>��THpn���kuб�K/��v&����r�ˆ��
�׊�1���v��:K@�9�&ۮ�=z9����Z��(N��O������7~5�� ���OI�-->�,8��$�H���b�s�0KcY*D�+�3�F�!.0�4̈z�����sF��j�B��W��)$����#͜~r��A��" ����o��bۜ?>��*T���jǜrr���d�b�P/9Ռ6����{�Rr�5�鵻K�O��Wka����H$^�D!�׹�S�@8��Yt� ���(A�g�1��ֿ���������$</��C�걐�|%؏�������-�y��������x��^]��`\�l�[���HWdڗ^O�K�o��a�V�}�_*}]�N���ȷ��AX�v%�>3a�I,e��/��$e�����-��3HaXz�J�^t���,���s>+]�2ںjGb�Ŧ�1���Y6�d��kޑ�6��8� �J�����O��s� ��a�Iv�ǰ�\���u>Jɀ�:��T�� hs��,&�{�~�ƹ_�&��A5�!�cz��z"��\)vC��R��XlxVHYEB    1f50     9e0n޻dLy�$"�mO *��#�-[�m~�˕;�J�h	���mV(T-Rwg���n;���7��Сco�$��6"�Y~	ᕓ��1������~�b䗇]+�L�9�#��.5��Z�}<��'q��9	�����{�󨈁^��������
)t����@�- a2E��Y�!�YY-�:�3�gBsB�n���/Fp#d���g��v�ݒ���m�nn�����vCsV�`㕵��X#T!l�_̽�1�RӮ��A�}�e�֩���`���*䐱cK�Ȼ��"b5�H��`��+�,���8?w3+/��3uk�1oS���ùQ����%��a����Z@��{� ��;L,1�mU�FZ���_��(x!�U���tE(ٖ���\�1K�g�p�[
H�/h�hTZ����3���O�Pi�\��ݞ0�*���hԱ[ſ��k�i_�-�-�����\`X���x�0�|�y0v�᜴���7So߭y�!�ama_S����c[�xF�)�ʒZ�.&���r����aգ,�D��t5�W�&Λ"mNo`�h�����w��v�}�6? H�i�X�NFO�*`W�Ŗ�ҩ3��+�2���w����&L������؈ݭ+����'�`���XY��C�<�N.H��J��c^�mg��^7f���tNxi�$@�?Mt8���q�R@E'��4�K��~��}=D�4�[@���u_�9"��BȈ��$rL������:G�k�S������M2�c8Րs�R��e���<��=��̃�џ��>��+�l����sn,��Q��o�����\�� /W���V�.��kDT�=��
����B�j0�V`�feQ#޹2�����t��q��n��� ��>S߬_b�_8��Z&�lK��]�q�)֊�e[i�`PM.�`�d��@ l�GCι�3:����zq�7� �K�����[�L��#])m��n���>�����F+tG���m�m��pѲC���\է	M7}�<ʹ]���C�|��I}v�u��Ec��B �5�'~�%��>us��9��2]���9R@��u�G1����GW1����'����֘>��M'���uB���Y���"�R��Z`�����Q&k[6oȗֈЫ�$�/ۥ�p�0�4'�������9���L�P�WG���������D]�ҏ �!lK>�!���Q�ڤ�1��o��ĵ�H�'��ך��`]@��}Ի��~7�2�]�'��'��/C�,�o�(xߙ�����aߴ8҅K����p�v�ơ�O���y�0�y��}%�>�Y����!:<NL ��i_���Br�O7L/`tT�U�������ޖa����.r�B�#����|q�ck2~�D���V\��+�8�@�0^�p{%&�4�ʃ����8I�����^��/�88E�{5R`�B�)� �Xf�<^�]�)X�Y�>΂���8�`z�)���B�!�`
1-���dAXX�MVit�J�+�&�4��� �������I`Rc�n�7�wS��C ���)k+c��í_2�7��*�A�s��C ��+M����(ȓlw��+���$�LMgiRSJ������%�R��fr�����Wˡ�A̔74���?��_�6i�����c�7ݢ�Q��������֓����Dq�/�'�Gʼ&:)�FV�����'͑��'o���=\ь}�["���M�!S*ӥf�G�@���LZ&"D��T��׳^��9'[P4f�C���5N;�ٿ��k績}�Cߟ����:9|r��F��t�����;���ӿ{���fכl9*�8�VKџ�$����q����X),s��q�V�r�>�C�cH�e��ܢVR\Xc ��
1�j�փx��a�8���߼�҆�`�q��B�0@&��_{R�.�Utx� |��|��>m��(X_�)~� G�c��/+�W�b��.i�/����3��S�L�\��|p�pk���)Gi�KΠέ[_�hCa�[���N��S4���l�	䤤�^�_5m��G�<���e���!�ą���&t��A�jЛ��-A�Gǚ� L�(�ܼ����Yu�����p����'�G��1pb����}Q����� �5k�s������T���sf!��!.���fV-�8�I~��`�-��4��0��c��U��+n:M�r$z����7���h�P�aO����H�.�l[�����5����C��G�lZ;yXT��6�#pJ�eaK��inw��mI�JHV�0��]�~d��!��W0I/��� �V�p����#�|uB%��c� ��~�4]G�pș
F��UNedչ��\ػ8D�}�t`�p��@�#��'+X������%U5 6쑨�[��৛s{�<�мoR��~~����҉2'�(P�q$`sh�
�p����B��;�#�}�g�p���X�n{�O�=>*?��-쒊