XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��WQ�@�X˹d߅�2��hS�ם�M�Fr���?��^�-4v͋* i�r�0@j��u���$>��
�KW����N~����h%4h&��E/ps�`�U�n;1�5���t��������>�qrU*l�)���c������'G�nu*�1���{�i���Et�G�����'�0n�5�t�V������͚�g ���s!��]V1v[R�G��R�����R�l�Z<����9R��c�!�/�g���Rp
�`�Z<xo���4C|4���8��"�4�[1^�Gο~�D����9_Oɑ��a6>�J�hB�2���
2XĞ׾��PJQ�$z�l���I�Q�|�r�a��+���(�X���m�m��X��阹�ԀѤ�a�j�ۧR��k��7��(Y�J�7��'�S��/�
�U6��*M��̀�02{��Jl%���`a�YTu3#��j�����B2�,,<_R:d�+�	� b�@Lp8zhM����_�J�2E`6ݞ�K�*���.����y���tb�jU�3͇X4`x��zQK�{8���2-�qM�AZ��6Z�y�بf�6�L<���/���P�D�)�i������@L�;�G0�<�Ř=�ǉFT�a����m���.��X~�R�7̙�M���Q��U�z:OE���2���ۚ�?���+�n�9�ݵ�N.�<�)��^�#p�4.O&���x/*QI���$\�5fr��`�,��P #��8�X�)�YXlxVHYEB    a04c    1c60�vs���5d̗&R,ͮ���{sP��j/L���e�đ��E$�_PzQ�jE�p)l�mYk�9�M�v_M�蟭������^l�����7�]��qV��^�N�k'�Z�r���#㓾�1�9:y��LVR�s������Kb$����G�\=OW����P7�����MϿ���X��&�,eb��7;�%�Iy����`�cPH��������t�|���~�~ЇV�X����vD�5>�}n���x�Y��=���/Ј�Ui�����	,� �
yH~�x�A�r:�S���i{��3��s�[���{��xs�DG��פL����^��#&��~�d&����nx���}Re��PX(O6��p<�Ȧ�<`��nv��a�>.VY'�d�gP��ǎ[����ՓvZ`3Ę�P9o�\́�l/m�d,�3
��DM���#�<�YNl�@a�*�CQ���v�i�6~�i1��^M&>��bU������V}�4r�����t �����ߓ�8��ŋ'�#qٱ�2��np_a�>� �,e(�B��B�c:X��>��!:�spK�������-�ش~����:���<��u���@K�2�͡���A�;�H�Bΰ]�:8\cY撫8����?F�����C��O�`bf�Xv-u(�!�"���8���T�$�>��:gywes��S�K�s�>s2�~޺�>���W^�"��8C.�?&���ųp���Y���\�|�ӝ�� =mt��A1�z�} U�ވ@�갗�6VX�j �gi�I���� �����1|Q�n､`��$Q�C����E������9q� S-���_M����>;v�]V�����ffd�ʆ,ȨB���I<:k,��JƗX)��ً�� �{��T_q%�����Q/&K����b��b�5L��{Y?ɕvߏ�ټx�x�I�V������N�0�BuX�-��� ���Ia��0&��������>�my�f� �ͷ�(\��	�S��m���Ǚ
���xd0��Q�k�ٽ�)�ĳS1U|n���5/���{IE���n&U�t ��ճ����&ȶ WU
�d�.I���� (�d��+���V�G�hΤ�U��Z��ü�֩vӣ�'�������o��3��_c?�Lt��w�M���o�Γ�h�Y�ʷ��h�r�-=V�tH5��*+��x�xfq��ߚ�ը=����V����dR��۞U,�i�i��NN��c�h{q�>�0����`$�ل( 8[�+�,����"���%��9�u�w?�&z8eU[�c:H��ھ��{գ�;|�L����"�ֆ������8�Z���IC�x�4h��-�[��7����=U T$�*U��| up��39����h�s=���+Gs�뗯u���l�1�KTV����0��L���B��|b�>���O��ɽg&�L$�E�(�^tX=I<H�}(��"�?B�>����SF�q�c�H��q=
�IK��=]�փr%��c3C�����]�O�$"�J`�CN�e��x"G�㾪CQ�����mZt����ؚyC�n�X���xQ��o՜F9��	�H�݄�}A�V�I�K&�=HHȗmަX�.w$k��/�)ˌ�9�߭�w\��/�,�4�*��Q |5�LIۻ�Rq���j�z�g�i�$���a�I{�]ή� �&t�7A���ҶQpƛ�NM����'_���?���7�u�NK�SvU_���Ӹ�u�� �0��*�ߌk�g�̀��J��6����]�c��~Ѿ�l3�B�҂p�+Vߢ�[�J�����ڪ�c�ftE@]�mc}�g`m���J�Q3w�C� x-d@@��FepD�a	^v|4�hĨ��`a���^���*@Zz*v
�t���$H"	vLN���sh����)իܿG��V�=��I8�Bj�<A�R���?Xj�C��n:X�W��AiF1�-�ύS�����ȟ^�)���]1�}'���K���<!,)Y�� N�C�kÑD����(t!�v��ҖDJ�	���b\�N���i�kъ�:/F�NsZ��4E;ķXHf�y\����{���W9|]8c�=0��s"2�~�>ڹ;�8�ѥӾs�;l���d��L\�G�	]�?�\c�>:p��8	�AV��΅K�ʹ찯<I��a�P��{��":���N�F�z>E)0�ی�o5�^�h	j�U?�_�>� &�v�E-��='^���k�;�.9�E�O5Mk����+9E䓩�o���/�`9�hk��;��#l�`m�t[ۇ��o��w+>X�l��]\�2b����[�?B�����u6H)�95v+"<�x�z����Y�I6j�ގ����sp�{m�����%�}���c0��m��
�jx;��.��੠o�C��wάi�i�}?畅�/�^�J��sv*D�x8Ͷy��8*�x��O�4��ӓ���]�"��ڥB�q:�4t�j-�� Af�y����z�K�X�F����Pz�1^\��	�"����v#�b�n���h�l����@(o&�է���RX�O]��uQ3z�{�R���8����F5Sw/gv�
��6�43Ew�T���8�櫿;~ۓKM��Ti/��3�4��'���+Yh���38�E�#yF��_X�;pM�����m�^�ڱ5�V� ��D�2T�s8��OQ�eKkN�=�ɷ!�D����G�Q�UԺl�`��&+%r1��Q*�8h�®�Z1x���R�?����V�l؈�P9U���\����%���	g%0��3:�B�%����M�	&�T��<��<:ۤ��l%�ͤ_�P�D�B�_��9�٢�F�;��c�L }��f�b\�"�q�s
L]�P�p">��YPcS�Ј�H�
s"��!Բ?W'l�(�A�o�y�oP)!�]�Yp�)ЈO��Y��r��8�.�EI�=dta��BU��2�{��~�y�ɬ�4���b��=<�����g������إ���� ����RmM��jn��Ϡ�!�Z����7BkM���yU3Π���qT��#d���<M��xf�z,�老D�S��I� ����2�6�S�m�>&&Maw�Go��\���pSOC��~"~�$�O�Dg�	* H�k#g�k�ui\1aD,IRM�'�f�L�z<W���G���銠k��ΜHd�� |#�%�X��ta�����EQ��l
�vD���cv��@&u7R{p����]ur/`��~&{�DU��jWT�-��a����b�S5to���N�b��nz���l��,�/���R���R7nM�1$f�CoF`��U��/)u-@wTHї�qź�~��dqD���/�QA��hG�U
�؜�a�#���m�&C����7�ok>�v���ȒP���J�i��\�|�C�zg�E�����j���Rcs_w��qe
%U젹���L~�ؗ���s+P�E1�Ay�T��_Ls��K�ˀ�M�O*ܙ@���\:e%�(�����(`9 ��b��DL�M@5��k���M��#PA������������L��DG�[��B��8I��R|G^c�UT�O�Y�Wbx�2�������Qՠ�]O(���_�@(X�����U�V�Ur� V�n)?�$*�N���}O^�}��n<��<�-RHA_^#ا�5��Yt��0j�1O�=�45�J��g9�����pA���f�����hND[�7�݆
�I���Ίg��������>�1rf�V��Ox�VѾrqL�`}-:��g� Ƥӛ!y�Na�7�Cʃ|&V���$���*����_1�wcm75�\͛�QS��>lN�NQ��Q/nA�	t�bw�A6+G�89m���2�7�uE�s�>.�����烙%{i��7�YTn��]�Vc�m��X��?q Yt�$6B���͢vD��J!�ze��&r�)�MUR�U�o	#T5�8��6���%��HZ1^��n�kW���jtkwVIH�=v.&y� �ܗړL�-��;��S�ʾ�$�J�k|`~4���%��b%�\����*�� .�b�~�)��A�B�riZD�� ��Ҕ�e���BG#X6�D�z��c��	�����;kA�[v��	�v��"Ua��&��������į��g#ڥ�~w)ǟ�f�%^�U?�84�Uլ�}��ɄdD� �'bf���^ew9��P�Gez1�y�Y��[�c�g�4�U����`�Nuf�.ǯ`1;�����n
��ٯW��-.bF<��wi�7����
 n�Q)a��N�ˮz'lO�l/�Y4?{gv9����h8IhϹG��K�S��������}8Hv1�\C�4T�v��i9�����2��80��I+��x�1������R]��
!�F?�x�+�?���{֖�ld*�};�d$X���@7R��c����!*���`�d�)�+G�_p����nyE?fj��r�x.�q���X��'�s�{y��\;�>�ޢ,�hq��uwn���Ͻ�Uu��q���|�i��A�4�;yc�89�y3�7&��̥�����K[���{{�%��Ћ����U��&���I���*n��i}��tE~ޚ��4��=hk��s����O�m�rg��H�O�'���ftG3��M.9W����bO�f��P��#�u qp�p�o�qL�B[�����B�0��5�c�f.E�6��=1��<�[���~F<L-h3�e��B\�ї�I�	c3�ِ7�OjV��i�5B.�g"�톮�����6�	ެva,��#	OM�u�n?��Pw�/U��{׳Ǵ��p�����l@R�Mg���~�50bf$)_�#����^��B��"��@�@��m�ȷ�
�d�\��)�	S�|(8�j'��n.���M��qCL���5�vZ�
�de�5��E�N��5�?ww��wW���V�OW���=T��xy�F�fO:���V��h��=��>�-��ʬNaDv��[ ,�+
�C�#r�V����(R�O��	K8�����A�+��d��Շ�P�ڶ}[���
3	m�`X��	j�t�2V�S4 +1�R�>F3G4��"s[,���w��`�yb�!��q�������'̘���g7T��m��93G� Q���������&[�ԡ@�m�%�)��]=,@r~x]*&�s��RQ�F�W9�Q�8QE��!SA@�퉔T�RKA<v7%(�5o�g�7��d+��Q^���j�E�G��%i/-)�ZXb��C�4�m����d���"���ɟ�GNآݮ`{4���G�"��|��Rؿ_��3�ݍ{�6VM
�~�*]f��t,�5��z�Ϲ�p�b;O�$���0���@�d�_e�<��c��(q>��[�} ,)��������]%�TG����7����L��+�N?[K�Xb
ځ�WlT���2��DF�{�����2#�ђ�����|U��m�$��r*��XR�4�:�xXy'�Q��LvY���%Gw��S0�0�n�[,F�.����`m�ݧ���S� �m�t�Yb ��]����C?��pq��=�8�#Y�b5��;��O��/vl��ǰ{�c|�4~uM���"��h�Ӹ̯�řX�o����&����b�
����Av��6��n[Q�z�ԑ� ��&�n�ڝ�1P����zU��q/���sٮ� �T:��)\�� L�.M��y���t��+��K�Pe�����xuq��s3&���5ٙ�yge;�)�k
+ �� ���Xav�e5�.����H ƏǦ��6���3�d(���m#%ւ� � ��^E7Y$_
?��Ð]�q�<���M�8�/?� ,���1H�(���3NW ��H�dWR��I���������k�;�N(p�w��S맱⦎l�~�mL�:�Zn�E'8������ ���K�F/����Hͬ�y{��D(�Y��[Δ����l���|������j;��\^>�g��ђ��Ʒ��8�i������1��r�������T�'!�ͅ�^�O�Y;f�N L����]!w����A$3�B��7.�Wƞ�&M�.Zw�ǔ�U$	l
��c7j0�QDm��y��3��^�l�qx>F���[bb�V�C H6ׇ��
�N�<��<f����X�[Ee���{�QVP��1F֞x�G�۝A�B5 �}�"���md�L
#{�@����-�DG/��{0n����<@C/6�z�Z�W��^'R�4t��@Zw�+�Ӆ��|9� q!ݱ�K3h����)f�3sb@��[��{}i�@n��'(�
;�j3'ǩ�}EJ�/�>�7��6���CH����棭 vr%"�Ŷ?�ϱ]�̭z��瀳ҫSX`�
p���{\&�o�@��sdE��v@Z�\I�+_��qw�^�F�M*�'��u&=��*��F�\m��W[5K?��j�3����x����v:5+ߌ���K�iqu��g�3�C�-z��ސօ�4c@]KZ��z�$����"�������r8n*r z�,4�jD{\NY��ÉA���V �R]U�5t���~u�o�����i���?��4Ȣ��@��˫}О{<��V~Q/NR��
b{ɿʰH�g�2��b�fT���0�ڞz��dk|($���M�ʰn[�m_s�tr�v�	��"��s�B���D������V�E��gs�'��Ĥf{A��o�h�z
RaW��:�@�MmE�H��0�bO�<}Cg=��o0�`w���-gA��^F͓E�)�;��?I>�ma��/p�|KP,��#9�:�e��F��r��PO?�{��:���������=. �ٙ�ԟ�@�>M���,�Ip�}�lCg��b��Նx�J��/T+�'�i����Ɓwsy�,�^����0���� ������o ����F?��:��f�I킕FXZ�T�c� �p�D=�$�e�O�0�y(]����R��<��;`м�	G0�		����{���g�\�G�����n�b�x�B��\���|[N��r