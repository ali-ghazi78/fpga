XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��z ��f��W&���7j~P�j��ċ��'nWb�VL;���@o����p\��|WQ��nbݲDܞ}��ErKFr��`q�S����P\3H,ڢQ��4t�8b�%ښ�O_�����K|���$D&.]iOk�MC*-�\�������A������"p�x�*a��I��)n,�i�N�����a�CR�4AFa�n<X��9�~�����s�0C��� :��u]����Vk,9��P�
ޅ�ǘ�n`���z�����W#�y�[�W~J��Tn�ʔV�ʨ7���O��zb���ϖ�TWܗ�d��k���������$�Q>��숡tQu[:���̈4�7��G&��y�t|?�Xj��K$����ɐ����o#��ʀ�fN#�|(�X�� [�B:��n��2���7��m�cFG/���$�	�����H� ��i��Cڶo�0�o��D���K��k��$�6_ɏnw(	�tU���&#ޚ�f$��:~� L�Z߮��<��OTw�r$�-T�q!���74�e�HuE�nz9�����A?�k��.���>���]�v}:���lΞV&9��.�V�����o"w��;����\�e���"�"�F�#���Z����=]��-�n�i�H�s��"ȁG!�`�%Y�b�U��#O�8@q�*#q�����|�2E�����M�^U񃻎ҳ�f$������r�������n�q�;���0s@�j�"[oN�Չ=$I�W8GX�AD�SB\��lXlxVHYEB    1351     780`eƶJ����2e"-0(�R��	r�E��Y����q<�%��� ��dB�bY.����֮Ӄ�{�%���t��G�Wϵ�>�#�p�gs�p�nz�c*|}��|�.����珉xkf*�_��}��� \^��Hz�����_�W=�_�.���[_T�%	��y��D�m]7^�j�ey���Yu��Q�	h�����C(��*@1�^���+!E�r��:{�gEC�d�9�ܾC�7:�ly�g.B�x߮�[� ؝�`;Vd]�l ��Z��N��;q�>�+Հ8�[(��h�t!̙�<���-ɺ�Zn��nyh�I%��\*|��,Qh��$�-���a��y�s��,%bhc�b�!s2�l�L�t�!,wz�?����<����izZ��dP� ��?��HEV��i�d�
�r��]=��D	�%*O�C>�����̥Z)'<$�O�2��������$yyI!�|:h!�)�`��?� �ų=�	�b"&S,w5!�7�ң����`1?$h��:�x�Ji �n� �!�mt���#cW��D�ÀH׳�v�J������\�4��\��m>JQ�C㴐�k��P�>�S]��P�NPⶰ���\��Z+���M�s�:�7G�䆭�qh�V,���g�)}�gb��g�|�	0��*��[�SU��1���+^,�i ɰ���_N� ,�$��A�/ͳ�,��c[7v�H��C8]�O���(�S�,h����{�1a���4�^"?��Q]��d�K+��_�w�q�����<O�	l��T���Hѫ��j ,�
g�f�{��F @�iT�m@7yj��iɼ�!�"�Ɵ�q�>��.�tU;< �����>��_�I�z��� �����w��5{[ul�<MM�Oߧ���f0�4�#`�t��s�F](=IG�^���s}k̘��i��_Բ�%�5���)��?ݸV��TS���/�5�����%�J���b������w �Oѩ�eVc�j-x�zl^�hoa��P7&z�+)3�KR��!��~Ŭ�=f��������IY`����K]�. ������G�z��2%7�\�`�L���v3�"@!���-$JC�6�E��ͮU�70���A�TD����*��V?[��7n�,a�g���$L�ؾ1�f]X� �����mR+�WY[>>�Y�M��]g�M�����(�ԠxmK�y]�Lo�����/�dov�~	���;�Mμ!����#Ltu2�o)%
���1#��W���YYX����3�m�d,����<�?�2hvMp���A��Z~�.�4x�é,�pc �>I�~Mq�G�*�ro?I����"��M�i맧3b�ՠ���ۤ�y�������
����-���ǹ�X3"�JI��)��d&w&C�P�%����H��q��<�eP� b-�I"\�b��ra�h�/�#�|����Y�w]���2	삔C.�ƕ��hr\�1��������7X�ݎ��	�S|X_���� (hi��I@"BȪ�*/�C1�a{},�u\��RAM1�c�rV�����N����r�{��O�U�ڊ��v�Q��%5�F�%V]�"؝��۞QP�$K2RzY�o�/ۈ�-�"ViN��;��R�B�L�'<� ;��;��S�֝�(�J"��03�?K\ �g���L�¸�>t�O�]t/�U�9�j�S��T;���0T畯O�����~��� �j�2/��g�E���K�ù�K*����'�?᫦�A!{Q�"��.,z�W����a�Py�[5T'�wT�q��ܔ���g��H?��#�+��a#$SEe���#�	qݯH_4�GR	����>iB�2�z�U�QN��c�%S}>8�ј���瓝@ɥηjf�