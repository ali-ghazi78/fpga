XlxV65EB    eee4    2910��l���a�GD���JO×B�,V�ɺ��]����-�hQ�R�%}դ�I�Z�v��ZqF�81=i���.P�1~��|D���t�?�2�k�������h�g�~' ����yv�g5��ݚB�#�6�qi�o�A����ҕޠ��46�h���"��#���j�ìgԉ�	A�U��X���,�����c�ƽ�{��"/�V{=�gU��w�����:@�E�ѫ�P�vL���I��� {]����P��6#yF=��$�@�a
5�3�3��a�5rЩ[0A��Bi$���V�<D]��Bt"�J �4'�j�	���F���`-�p{� �( ��:����$�8�e4�uMc�����?N�#�ؗ`&��*�?��.ptcx����6�Ne'r���_\kw,�۟=nel�@uA��!�Qv��&.�:j8��b��'���_��|N����b�%��+{���$X�	�����X��C���3&�>(��=��o:I�vz��M\7��&�%#V�:SЂ�i\�6q�xB��4.2�v�p���UG��@AT�r$ ��i�0:I]ϯ��#��4vjDbW:���|u�!r�n�Z����j�])>��`i��Rr2���z�����qa���71���<	QN��ү���k�L�}"�v���EM��KRү^LmK�	��`����p�-tZ(p��c�K,�x:�������,�0&^�Ib"�^�j	�۷���֮N�-4���Jo���i6u�-�&���	��y3��.Qj�(��'l��^���\MJ.wφ��� �Z�i���s�j|��x>��d�̱h��� >����m��S�Q���{����LԂ��d�i�� ��}gы*ww�z�%\�d��E	�^����cr�*(h��:������A��c�$:A��e���Q"��-�h2mgX�r� ���04"�8�������\�S������x�d��1����a���Oڃ�F@�t�>��l�B�Z�:���ew���)�v��l>�NI�ad�)z�a*� ���D02���Q�5����oh�xA� U
�?�!*L�a �c%�d`�]y*�����W���q��my�Q�5�B�z�;�z�W^�>�?豽Hp��:Е�7[c�'�[�;���g�M;޽U\�u��̿��I��vˁY�y�17>{�u��1D�q���0�㪑�*l��+�z�\*����7�p 63��3��f�'n��O��@%�	,��PVD<P�����ݴ]H����d^[r�I4�K���x��j�v�� q8ͱ����[�~m�����iUY�M��%�M^����gjd�{
�D�=��ms�*�h1�9��2~52%ռ�����{�a�#�j��/X��Ԭ��Bw�o����"�j�����Q��ԲL��������L�ZR3q�Cv ������ӵ�|�䈎��N�a��5F�;����郷
[������k�h#Cd;����6y��H7?j�6x��<Q�H�mq����X��ف�+X�ٲ_H���?���`,�6�Y/���@���o��	/�)��Y]�B��b�X!�C��e�*�z�:��R���Odgd�\ppfI���RF�Z��i�M�d+�F��S�g6*C@>���&Gcw_��}�F��ƅ�����ǝ�:JmW��b��5F���I�xp�H���N���[�0VwP5��������@N��=��̸
��_�?�ʨ��)�U���~p��oQ�9A&Q�9nFT�H����w���6���6>�-d>[j���bd��H��@ *��2��-ț�M���8�E�W@���2*-Ekd��c��+�L!�u�qH�����$Ѱ�u͖;�m�P���N���0.��Zsn��Ѣp�z�`)�Ý�8���Eng�~�]��Rx���x*߆��~�+?8��(��y�%͞���I�V߃=� f��4LL&<#�2����wo�-�	hJ��fɪh<�2-2))LZB��#���R� )t<��2��D�ຬh�/�F��fޗ��u����	V]B~T+���yJ�@�F�B�8��2�yu���h���d��c֦�!��[�D����y ��b���lYHϴ�<*���~&����� \�� RB 4d�n/q���3yv�xh���_�W�7�<v����
�Y��R, ��끫�?ш�R��Âڀ��7�!K��_�H~M*�}�c:���z��YOpͨ���p%��FN�y�p�q�'b��
�w�k�޷B��9��E_[���ǳ��#t����0�с�9X�9!^?��Ϙ��)�)JHr����S���/��� ���Yc���;Yo0Un�ݾ9]��E�	�Kv�R����L��4�*[������b��@��V.�0D���ʂw�@0e	E�U;^������e�ɬi�
�ЉJ%C\cKdx&�r��D�>+���a�'�+�m�@Sx$^b1�L'���Lh��u��U���c���xjNF���A@8��0�l������<�:�6����9�,�b0
ڑ�
.���H	=!'�4����.�������3B���h��4���3r�h;e��Zkf�_p(qpN�'��<�������vk�{��$کU]<���J^La��˻D�jk���
���נ!TUo���Kɦ���d��V��̐��9;_�0U���7Av)�au��U�AL�5�cԒwԏw�7���*q�޺�&�۔�Ā����ʍW�mhbN�>e܃m������R�B�;ȠH\��z�<�Jz��V���1[�?*�wGb)��`^�;�x��U���5Q�c�/`�CH2�2yO5�����g�[>
8�R��'F�t}�V��~���^_ ���u�������v�o��|E�[�3F�����I�Q��)�{�KKO�i��7�L�����6"G�>A�5���W������Ke�w��~�?f�u)š�f@z���ĥ��P�U����rw��٩[�*͎:�\h]���� nxq��K�ƞJS�fP��H���Zv�V�ԁ�#f�+xd��pQſ�Ek=�r ���cq�2�j��=�C,��P�E:3��W*)�4����ߧ_C��?�É��菠���v��Љ�%^���kƜv�zE�3l�qJ�e�/�V�����%��ˀt�y	��ʁ�?�u�._�(&х�]���/��!��+��;Kw��k�*p;+�HI����)�z�Ph�a�YTg�$��A�|���$-Z�\5��e�WHt��P�kTDB	�F�TNO-<�J���%�7񛏭u ��t?��Ԑ$,�p!��^"hP4����.�%AV�Zq��$\xm�:�<+Ӯg<r`~r�]rC�D�=�f>tk�͐ȸ�_��a��/��T\q�N�ZQ�u��ItLS��*���]���_��P��t��J>��0��"/}ϟf����~N�u=}>
7�XA"'�i�xԇ!��"�ek��E�i<�A�V���AҢ\xsW�.)¢5���T)=#�w� �p4XR5�ɹ���s�l��eqb����w'�"?���"�)�u"�b�y��[���G���{�3�x��U����D�~��V��Q���=��~vk����yJ1Q�� �JI���䒇[��^�0��|)�� ��+@�>[���"�?��K=��/u䃧���C�������|�����E)��ԕҲ'U2l��?9����:���g�ӡ�H��i2dIE"�
k)|j��/?-Gx��Z�1�*M|��|��!e=�;�E|��/��藢|^) �+����a��8���QF��9���O��1��7���ޜ�jZ+e��#)��fa"�0�j	9p��V������oT��m���o:��ΫO&R]Q�02���s���j~���P�BK}���R
,�Y7��|�5M����;~*�R��T���f2�ɢ����Gb��7k�c���6���Y����H��T5���x��S�x��1_�P�*C?ﻕ}[�U�~�?Y(����rNw'V4�xp3���"V����IO2�t'�M�6U�xy9�<�sk�XЂ%����������%jGP	^��T�E{�DNb�!�M*Í	п/犷���HJbx2T@HT��x�Y�+��*��(��8��}��]��_��2:Բ#�"��@���\/1p��&���Ix�<�r*F��l8���]sOCxN��T6�k`���)珻���Gu1`��>���]Ў�)����V�Y�"mu�F'�s���	 ��&K��T����v:��A�!�5���Y\�.|�f�6z�2���������e,SL@��vF7g��"x���꙰B� Q�2~b��0^��Y�)	i8R��7S�K̓�+@�v��ďI����J�Ѧ�z�j����3��������_i�����3����A�l���sR;󼺹B�
VA/�ف�9��$�/%��!v�xv�A��F,���كѱoSQ�+{\(�ӭY20&�:yXⰡZ|�X��ම�I/��8�5Qe}垲,���ܹ�sd����.���2�u�a]�m�ǂi�]�Dd���<�;l�	�i�Ӈ8��R	炖�ܨԬ����5�e@ݶG�ϵh��M���/C�l7I� ��E^�b�\��W�����y��##?������5��^̀�x�m�r���0Fs�4����B�HV�Ys:����L��O�� }O����;�X��4�G � c�0!��1׷Ex��]�TX�5
(NdYR�P�ߑ����1��������i��i�q�^!�`���N)�ʃ~k���!(��u�b����O��&C�<ZF�����<5� �88���e�!�7��h��O2��4'_F�z���"g�k�-�qSg���-3� KP���>�d5�>�a5�;0k���N����E��g��˰8H:S{��kEn�o�\ҧ��k .A.(Zz3OwL�"UIs��9*����#���O%`��%!!1�o�l5�.�pNh�862X�&W-k���kO�-9��R0TVt��C���n\s�Z��c@ޯ��p��Pxd\��eF�͟���2AOS�����S�S߀\5b�^�v(�t�-�<�j%��q��u}��|m���������p'� ��7r�����>��hNTrcq�6�S�Q��28�R]�VK�+s��P����l2�vDXb/; -���g-9��������n8���
 FԺ@lx�j�gޛ7��t���V�ߛ��f҆#B��vw��#:w�[�f�!ݤ�K ��N��?����#Ein �]��\V�Zv�|46����WρJ߇\B�ޮ�"#t�|h0�A���o�(�W�p�4����c�ar�s�~���Po��1|�������j�KE�BJ��,����*Y�C��Jo-���TYbe� ����Î� ��R`C�l����J��{\�d��j؜��~�!�� Xm�	����
h^`���ªp0�����8f+Oy}:�.�@,�sK�67�>8����pʚ��n	\M)����۪}��?E��!�G;S�pj���481D8_��؜�=Y�v�N�v	�}��W i��1��☞/��� ��������4��+�zAt{$P�u�p	�X,�/�͏��F!����.��i��j܀��gk�g5tYk��r���,�<�_� �?�G�y�����Î�8h\�~��M�Y���K�ܠ�|���1���4�P��[�
w�ۼgL��ȿ�iʣ�:�(���jP��C����p�7�����tiL}�mR�Pd���|vϦ��Ja� ���1~��[��͵�p�&��=�������*���{ZX�4�ƅc�Q�,�r��4���L���cv���;Cj�l/	/��6۴���z���%��-Z@w�$K����1Ok'	�S�.y��~ �3v=���S`�Wj��,-3���v��;�K����g#�ceN�|��	nnG�n�P�d���	�b:O����3���xhI�@��,Zui�3BU�̧��f���>;�Ez�`��LwV-O�<Ay
+��%�Q(͖���z�e���ϴ�����dX�]HoL\���!�ϘK8l�gY�����'r����:�j� o*切�lVn��#�(��S!��#�N�8T^D�1��'����7`ғ�0&�KS�@o�c{7���'(��߅���(ݍ�_��G�?��� ��'�b@W�}��ӯRY�e+���*n��4�f3am�ǽ�l�ѶަɄn�9@
c�7e2�f#��D�`��b�Ya��I�W�h^��~8�O�<�����K@)��ǥ��,sU"��B}x�#�W	�m�"[�;����4�LK�M��y���a����G�C�K���Gg�7u��W �(xRؔ�uO4���P�t����݂�|�����5]�&?x�nB�\�O {������{j�����Ө��e_勦�l�Y���gC�_�5r��������Eqk��C���:I�s�*'>ӂWU~}{c'[��Ñ�3�4�:�e̰
1ж����� FdCH��d�)� �/�ʶ���LBl��7����W�[{�mu���o��u=ۘ ��$�S4��&gZ�0���H}��cba^�Ҹ�
i��u���<��$IH���~Q���8Q;YYrKg��up�s�T1��#13��x�g`B`[|�����Yo7�KX�	Zk:`�k�j3r_�@��"��N��?��|.c�Z�y��N����?F��6��C�`nF#����_!�b-֧ѓ"��Ĵ�f��<EAL}qIl����+e��Xf���7_�v��.n���:R;� ,���Wg�:�#��W?ڮb����%=� D� LLAoUz�|���ҴZ���/��sl�e!)w��j�nq�]�H���q̀��{��>��l0�����[APh����0���	�u ��X�R�|1G�j�WK������	V*�3Lc�]M ���ͺF�YX��)���RH���ĕv�N|��\��Ը�����"�'qL21����O��r�$�O�ً�_&��G#;X)zUs\a�b���e�	�=�7�:��6���BH������-��<;u����J�Un����1���B�:y�:��!>����(5���$����4�| �Z���;��/SyJ���6GB�����Q1w��lzK�0��N�ى+�,u��*CՖ��Ƅ��4��6�P��'{l���g����֪j�8��2���{�:�cw֒�S��D'�DS�w����G6��f��+�����-�K�5����s��y70��b��������}N�U�@.�_�b2�2;�-������(�U��N�<x�B�z���wq�Oώh��2"�*�����Ì^qT������Z���c��7��r ݫ킮�{��\�Y^�WP��Ӹ�c��//��'l�4"Z.����O�xhg��i���.
�y�1ܧμA�j!�Q�k�C�K���}(������/�J[3θţQ��Þ��~8+v�Q�B7��hg�Lgl��΍)M1�]nM�Sk"K?Bm�pvD&��t`�E��8� z��Ȭ$��`2��&��}wG�lAQ����	v),��w�w�t{J�Y�:�z,�LN�h(C4z�����v`�Hk%�VK�=U,��h镡n��|������-l@���f��:�oY���FV�Ȁr����kU~��������v��XB�Sh���`p�"l?��z�CV�I��K��\�O��!#��[���x�7�fb������fm��0�^�F�3����J����Q�s��~�JG+@��PtI����U:�g�l�˃3dJ�b=S�-��'�wo�X��7�a��RCL��nО�N�b+!� ����3�HB\~����U�H�(9�w�@$f<�=��ӰO�f����HAZ��!��S��2!L���/e�/;��a5GD^����tdE�uB�e�11��!��M89��$�����Yܐ>+wiR�gI(��k��T"�Գ��	?.��H�8iH�;"������}5��v��i�&��ΫPp6�tdsabX���(��ר_����L@��j������ZR$��Nb�� ١���'
�c�~[<[k��$���fZ�f��H�j�� ���ԛ�����0H$I2��C�@�ˉy�i`�8�SEStyP�l������v�u���W�`Π�e��"|�W�*��S����\mr5Z��z�Β��9!�8���s�%X'�aO�k(˶��[1F��$͆�e�6��JeW���pC�[��U��������ír=�&==yh8͹#��T�[�dZz�ʥ.�F�.�l�m�Z��*gF�gF�%�J�f砗��|��_ ��8�����'��Oq9d"��\e��VK������vN�W wZ���=-�B�"I" Q%ߕ@�p)�z�E4�w��M�E+8k��N�,�/��\��;x݃�@leI�,c��`��8hJ�]0on�X�$S��r��F���Uٴ�F�{�54&�9�c�I�5�����O"�C��0` �/�<�(���:���c��n>tʦo�۩	�0[�5��G�V���ޛ@S�΀���� ���Z���*98`i!��W衐�~<���@���.�Z/�	'��F�������rG�@P���t����|~p6�g���[m6y�!3_8��M��F�YԢ���ydU(��&�hY��%inIn� DVf��t��0��V|X�]��,����\�; Y|���+S��p�9X1^s;��!�T_�a�+��嚾BgG	�TNOGD�W�:��Ata�ƌ��R?_��D~S���/2я���E��O��6�bξu��ßIױE���H�TC~�&6��'q���i�
��@�@U�=EWu�>g��K&���m:F(ݰ������������Pׂ���ʐ�u{����H�B�G�Ӷ0����co&� �f\�|O��&)������̑Q����{�� �>�!gn|{blg��db�w���wx�X���䛏�~��7����F�ҧ�^�E�f�H���F��t ��˿aM��兏��2+0k��
~>:��x���s��@q���t�w��/���;nn��k��UZ���qQġ�Id���t9��f� �1DG�,�1G�QoExe��BS~��ώ,��~5���V��L��	���S��{����G��z�z�􎂢f���+���mYW��J���q�R��/��>V�Y�\�f�����>� ,����N��YR~����ٴ��0p�����Q䮟2H_����������\�U�3���A�1t��!zm�k��~k��¨�$��ɱ�����G�]ԇP�{��S�����:$-�k�VC�@�D���ʋ�ㅎi{�3�k��o��	�Q�]n3$l��������L*t.��k�*��U�JH���o�cQQv
1tPIJX@�$[��[ڐ)x9�H�s��ZC����w�'���8ʨL��7�F:�p�ȳ%�����9y5��w[��'�����Bg���lv�y��[��]��V�&�Q�Q�*�m���󤚿�Dc�i�B�DHr�^o���!��Q�L���V%7kxw�8��>�n�b����S��V����+��o���>
yH���x��+8*�ͧE��p�v^*b��QTa͆�p*G9{\pe�a}^a��23B�j�ǉ-��.�B���}�o/�(����y#���J�����A���Q.���El1l��L5�=��9�H�Ҡ�߬y���qw��_n��_X�Wv��ҟl�pac&l2̙5�nٰy���b�z-]�m��MSܴ�� ��܌p¨��P�2��0����o߾��K6s.RZ�<�O�(*��׈�}
iw'P�)�����8��]�ho&�,E������2���'�A�S�%�i���<q[��D�j��S�:¬��:����h��q�R!��p�ٖ������6pLlƮ��<�{�$�B�8�p_�Dv�yIz���A��̟�c.6!�?b�j�v���-�H�Ƀ~�Z{Ḙ��+���8Z��g6�m�t^?b63yD�)1m����K�a�sa���ag��5�gK�m�1��y7�%]�B�h6`/���qc	���8���I���VN��e*x�eF�e�Q��\w�O�~�a�y