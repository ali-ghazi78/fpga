XlxV65EB    1350     780&ه��Q��O�Tڣ��\�?�;�cl ���8(��8�[�7���V�8���7Efw\�C����~
�2�i,�}/��Φ��b'�9\��2���2h��Y]��>�!猪#W�T��#���4��T�/�損���R�V4cXV�1U�_������5v��.�*Z/f��unJ�~k._�:�ȉ��q'�)��Jy�q}��-�N|��Thڔgg���|wթ����j�qaZV�w0uf~�{��l��?c(�����S߽�W�U��\��OXr��>N깟{�=w	vӲY�{07����
!y�&Ӝ�{0�x7A>]q�I*=g�&��?�������qa�P���a��3B�ch��F�?�d=�.���H7":P�cP`���;�w��r�3\=@��^|�*եT�Yt���R^k!�j8�Y݁�9��+կBj�5\�B_t�NC�8�÷�8�����<�a��~͍2��x�w�s�:wc\�^�Q���g��a��Y�2sD-D�)kYh�� u��hlj�7��P`��2�)�4�����O-�]��<�*g�4�^�ƪR�xq�W\�/ƌ@)�LZ�!~�N9�޶����aפ`��`Cp��}�@�1_b�}o6�eT���7�^K�Y�P���Td3<�n	�ٖ��Ԥ�3Ya�|�U+�͎&#�3Ḙ�w�s�UR�u|�MA�>'�y�X�VJ{y-2�H%�_.�@���j<����ˈv�s�D�tܞ���Vc)�w/��e�����t�+��t���{øH]�?Ȋ��<���Ĵ(��[��1��EX��*�>)7A���Z�6�V6�w�b��:�
}
�^��{Ũz8�C����g�}�srm��M��Y���?�q0l�	��a9��R�f�󓰔!������@3%W�j�0�a^�C#~'�|���2�z:G'Y�#����Gyu��i���u ����2�
.�/��@�ʍ/���ƴ!���F�/��!0B����*Z�|����^Ǌp�<�-�7s�ĘD�G-�>�@��� �4g�
�6��G�L[�og3�3qu.���EV�v�	Y�"M�Ef�Q6��}2u��]F�hL-S��^�}�LO�A�Q
�{��~�n9>��Z�Mq��1��	*yv��f��=��}���������zw����hUX%�>W����U-�B�H^V
��}�~�)���W:�Ge�C��g��k�H��K�mJܠ�[���b ��.���7Ɯ^_PL�״��C��h���E�@� ]�H\J1À�40ӿ��-�1���&F��#!F}E�rGX�(Z|V~y2R*�z�ϸ�0"yd��<R`���Z���=����q�I|�@J�zv���x�l��K�F�YN�s#��l;�c��.B".�ꋏCUv����Ǹ����`61��L�4���"����\S�Q���`]�;�	��������7<(��~q����	��H������Lh�Zɠ��䫹���#"0%N����{��S��]�GĆG� l�ɪ�t��#Έz*&�ߊݙ��ؙ1�h4�\0������9����0�����m�kU0XB�kZb!,m��,a�oo�Sɨs�}�Tk��]ʭ�<�"q�Vl!���[H�;� ��$=;����2W�t����޹�\�M�����HCi�o�Cx}1�M{���J'�����H~/BJ��q	y C�2�p�+(l�ug�D�P�cm"��A���-sS�`V��>Pڎ0_���~���j��G�'qK7����%@>x	�������ޚ�I�iK�a����"���R�3��偊/!y��\Q���ֶ="SY�	��uC� ,�x�>a;	����ݟ���*|4�p�NV��tC&ɋ��0����XDC:�o�)����1d